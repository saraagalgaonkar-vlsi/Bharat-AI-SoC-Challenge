

module yolo_backbone_accel
(
  input CLK,
  input RESETN,
  output reg irq,
  output reg [32-1:0] maxi_awaddr,
  output reg [8-1:0] maxi_awlen,
  output [3-1:0] maxi_awsize,
  output [2-1:0] maxi_awburst,
  output [1-1:0] maxi_awlock,
  output [4-1:0] maxi_awcache,
  output [3-1:0] maxi_awprot,
  output [4-1:0] maxi_awqos,
  output [2-1:0] maxi_awuser,
  output reg maxi_awvalid,
  input maxi_awready,
  output [32-1:0] maxi_wdata,
  output [4-1:0] maxi_wstrb,
  output maxi_wlast,
  output maxi_wvalid,
  input maxi_wready,
  input [2-1:0] maxi_bresp,
  input maxi_bvalid,
  output maxi_bready,
  output reg [32-1:0] maxi_araddr,
  output reg [8-1:0] maxi_arlen,
  output [3-1:0] maxi_arsize,
  output [2-1:0] maxi_arburst,
  output [1-1:0] maxi_arlock,
  output [4-1:0] maxi_arcache,
  output [3-1:0] maxi_arprot,
  output [4-1:0] maxi_arqos,
  output [2-1:0] maxi_aruser,
  output reg maxi_arvalid,
  input maxi_arready,
  input [32-1:0] maxi_rdata,
  input [2-1:0] maxi_rresp,
  input maxi_rlast,
  input maxi_rvalid,
  output maxi_rready,
  input [32-1:0] saxi_awaddr,
  input [4-1:0] saxi_awcache,
  input [3-1:0] saxi_awprot,
  input saxi_awvalid,
  output saxi_awready,
  input [32-1:0] saxi_wdata,
  input [4-1:0] saxi_wstrb,
  input saxi_wvalid,
  output saxi_wready,
  output [2-1:0] saxi_bresp,
  output reg saxi_bvalid,
  input saxi_bready,
  input [32-1:0] saxi_araddr,
  input [4-1:0] saxi_arcache,
  input [3-1:0] saxi_arprot,
  input saxi_arvalid,
  output saxi_arready,
  output reg [32-1:0] saxi_rdata,
  output [2-1:0] saxi_rresp,
  output reg saxi_rvalid,
  input saxi_rready
);

  wire RESETN_inv;
  assign RESETN_inv = !RESETN;
  wire RESETN_inv_buf;
  reg _RESETN_inv_1;
  reg _RESETN_inv_2;
  assign RESETN_inv_buf = _RESETN_inv_2;
  assign maxi_awsize = 2;
  assign maxi_awburst = 1;
  assign maxi_awlock = 0;
  assign maxi_awcache = 3;
  assign maxi_awprot = 0;
  assign maxi_awqos = 0;
  assign maxi_awuser = 0;
  reg [32-1:0] _maxi_wdata_sb_0;
  reg [4-1:0] _maxi_wstrb_sb_0;
  reg _maxi_wlast_sb_0;
  reg _maxi_wvalid_sb_0;
  wire _maxi_wready_sb_0;
  wire _sb_maxi_writedata_s_value_0;
  assign _sb_maxi_writedata_s_value_0 = _maxi_wlast_sb_0;
  wire [4-1:0] _sb_maxi_writedata_s_value_1;
  assign _sb_maxi_writedata_s_value_1 = _maxi_wstrb_sb_0;
  wire [32-1:0] _sb_maxi_writedata_s_value_2;
  assign _sb_maxi_writedata_s_value_2 = _maxi_wdata_sb_0;
  wire [37-1:0] _sb_maxi_writedata_s_data_3;
  assign _sb_maxi_writedata_s_data_3 = { _sb_maxi_writedata_s_value_0, _sb_maxi_writedata_s_value_1, _sb_maxi_writedata_s_value_2 };
  wire _sb_maxi_writedata_s_valid_4;
  assign _sb_maxi_writedata_s_valid_4 = _maxi_wvalid_sb_0;
  wire _sb_maxi_writedata_m_ready_5;
  assign _sb_maxi_writedata_m_ready_5 = maxi_wready;
  reg [37-1:0] _sb_maxi_writedata_data_6;
  reg _sb_maxi_writedata_valid_7;
  wire _sb_maxi_writedata_ready_8;
  reg [37-1:0] _sb_maxi_writedata_tmp_data_9;
  reg _sb_maxi_writedata_tmp_valid_10;
  wire [37-1:0] _sb_maxi_writedata_next_data_11;
  wire _sb_maxi_writedata_next_valid_12;
  assign _sb_maxi_writedata_ready_8 = !_sb_maxi_writedata_tmp_valid_10;
  assign _sb_maxi_writedata_next_data_11 = (_sb_maxi_writedata_tmp_valid_10)? _sb_maxi_writedata_tmp_data_9 : _sb_maxi_writedata_s_data_3;
  assign _sb_maxi_writedata_next_valid_12 = _sb_maxi_writedata_tmp_valid_10 || _sb_maxi_writedata_s_valid_4;
  wire _sb_maxi_writedata_m_value_13;
  assign _sb_maxi_writedata_m_value_13 = _sb_maxi_writedata_data_6[36:36];
  wire [4-1:0] _sb_maxi_writedata_m_value_14;
  assign _sb_maxi_writedata_m_value_14 = _sb_maxi_writedata_data_6[35:32];
  wire [32-1:0] _sb_maxi_writedata_m_value_15;
  assign _sb_maxi_writedata_m_value_15 = _sb_maxi_writedata_data_6[31:0];
  assign _maxi_wready_sb_0 = _sb_maxi_writedata_ready_8;
  assign maxi_wdata = _sb_maxi_writedata_m_value_15;
  assign maxi_wstrb = _sb_maxi_writedata_m_value_14;
  assign maxi_wlast = _sb_maxi_writedata_m_value_13;
  assign maxi_wvalid = _sb_maxi_writedata_valid_7;
  assign maxi_bready = 1;
  assign maxi_arsize = 2;
  assign maxi_arburst = 1;
  assign maxi_arlock = 0;
  assign maxi_arcache = 3;
  assign maxi_arprot = 0;
  assign maxi_arqos = 0;
  assign maxi_aruser = 0;
  wire [32-1:0] _maxi_rdata_sb_0;
  wire _maxi_rlast_sb_0;
  wire _maxi_rvalid_sb_0;
  wire _maxi_rready_sb_0;
  wire _sb_maxi_readdata_s_value_16;
  assign _sb_maxi_readdata_s_value_16 = maxi_rlast;
  wire [32-1:0] _sb_maxi_readdata_s_value_17;
  assign _sb_maxi_readdata_s_value_17 = maxi_rdata;
  wire [33-1:0] _sb_maxi_readdata_s_data_18;
  assign _sb_maxi_readdata_s_data_18 = { _sb_maxi_readdata_s_value_16, _sb_maxi_readdata_s_value_17 };
  wire _sb_maxi_readdata_s_valid_19;
  assign _sb_maxi_readdata_s_valid_19 = maxi_rvalid;
  wire _sb_maxi_readdata_m_ready_20;
  assign _sb_maxi_readdata_m_ready_20 = _maxi_rready_sb_0;
  reg [33-1:0] _sb_maxi_readdata_data_21;
  reg _sb_maxi_readdata_valid_22;
  wire _sb_maxi_readdata_ready_23;
  reg [33-1:0] _sb_maxi_readdata_tmp_data_24;
  reg _sb_maxi_readdata_tmp_valid_25;
  wire [33-1:0] _sb_maxi_readdata_next_data_26;
  wire _sb_maxi_readdata_next_valid_27;
  assign _sb_maxi_readdata_ready_23 = !_sb_maxi_readdata_tmp_valid_25;
  assign _sb_maxi_readdata_next_data_26 = (_sb_maxi_readdata_tmp_valid_25)? _sb_maxi_readdata_tmp_data_24 : _sb_maxi_readdata_s_data_18;
  assign _sb_maxi_readdata_next_valid_27 = _sb_maxi_readdata_tmp_valid_25 || _sb_maxi_readdata_s_valid_19;
  wire _sb_maxi_readdata_m_value_28;
  assign _sb_maxi_readdata_m_value_28 = _sb_maxi_readdata_data_21[32:32];
  wire [32-1:0] _sb_maxi_readdata_m_value_29;
  assign _sb_maxi_readdata_m_value_29 = _sb_maxi_readdata_data_21[31:0];
  assign _maxi_rdata_sb_0 = _sb_maxi_readdata_m_value_29;
  assign _maxi_rlast_sb_0 = _sb_maxi_readdata_m_value_28;
  assign _maxi_rvalid_sb_0 = _sb_maxi_readdata_valid_22;
  assign maxi_rready = _sb_maxi_readdata_ready_23;
  reg [3-1:0] _maxi_outstanding_wcount;
  wire _maxi_has_outstanding_write;
  assign _maxi_has_outstanding_write = (_maxi_outstanding_wcount > 0) || maxi_awvalid;
  reg _maxi_read_start;
  reg [8-1:0] _maxi_read_op_sel;
  reg [32-1:0] _maxi_read_global_addr;
  reg [33-1:0] _maxi_read_global_size;
  reg [32-1:0] _maxi_read_local_addr;
  reg [32-1:0] _maxi_read_local_stride;
  reg [33-1:0] _maxi_read_local_size;
  reg [32-1:0] _maxi_read_local_blocksize;
  wire _maxi_read_req_fifo_enq;
  wire [137-1:0] _maxi_read_req_fifo_wdata;
  wire _maxi_read_req_fifo_full;
  wire _maxi_read_req_fifo_almost_full;
  wire _maxi_read_req_fifo_deq;
  wire [137-1:0] _maxi_read_req_fifo_rdata;
  wire _maxi_read_req_fifo_empty;
  wire _maxi_read_req_fifo_almost_empty;

  _maxi_read_req_fifo
  inst__maxi_read_req_fifo
  (
    .CLK(CLK),
    .RST(RESETN_inv_buf),
    ._maxi_read_req_fifo_enq(_maxi_read_req_fifo_enq),
    ._maxi_read_req_fifo_wdata(_maxi_read_req_fifo_wdata),
    ._maxi_read_req_fifo_full(_maxi_read_req_fifo_full),
    ._maxi_read_req_fifo_almost_full(_maxi_read_req_fifo_almost_full),
    ._maxi_read_req_fifo_deq(_maxi_read_req_fifo_deq),
    ._maxi_read_req_fifo_rdata(_maxi_read_req_fifo_rdata),
    ._maxi_read_req_fifo_empty(_maxi_read_req_fifo_empty),
    ._maxi_read_req_fifo_almost_empty(_maxi_read_req_fifo_almost_empty)
  );

  reg [4-1:0] count__maxi_read_req_fifo;
  wire [8-1:0] _maxi_read_op_sel_fifo;
  wire [32-1:0] _maxi_read_local_addr_fifo;
  wire [32-1:0] _maxi_read_local_stride_fifo;
  wire [33-1:0] _maxi_read_local_size_fifo;
  wire [32-1:0] _maxi_read_local_blocksize_fifo;
  wire [8-1:0] unpack_read_req_op_sel_30;
  wire [32-1:0] unpack_read_req_local_addr_31;
  wire [32-1:0] unpack_read_req_local_stride_32;
  wire [33-1:0] unpack_read_req_local_size_33;
  wire [32-1:0] unpack_read_req_local_blocksize_34;
  assign unpack_read_req_op_sel_30 = _maxi_read_req_fifo_rdata[136:129];
  assign unpack_read_req_local_addr_31 = _maxi_read_req_fifo_rdata[128:97];
  assign unpack_read_req_local_stride_32 = _maxi_read_req_fifo_rdata[96:65];
  assign unpack_read_req_local_size_33 = _maxi_read_req_fifo_rdata[64:32];
  assign unpack_read_req_local_blocksize_34 = _maxi_read_req_fifo_rdata[31:0];
  assign _maxi_read_op_sel_fifo = unpack_read_req_op_sel_30;
  assign _maxi_read_local_addr_fifo = unpack_read_req_local_addr_31;
  assign _maxi_read_local_stride_fifo = unpack_read_req_local_stride_32;
  assign _maxi_read_local_size_fifo = unpack_read_req_local_size_33;
  assign _maxi_read_local_blocksize_fifo = unpack_read_req_local_blocksize_34;
  reg [8-1:0] _maxi_read_op_sel_buf;
  reg [32-1:0] _maxi_read_local_addr_buf;
  reg [32-1:0] _maxi_read_local_stride_buf;
  reg [33-1:0] _maxi_read_local_size_buf;
  reg [32-1:0] _maxi_read_local_blocksize_buf;
  reg _maxi_read_req_busy;
  reg _maxi_read_data_busy;
  wire _maxi_read_req_idle;
  wire _maxi_read_data_idle;
  wire _maxi_read_idle;
  assign _maxi_read_req_idle = !_maxi_read_start && !_maxi_read_req_busy;
  assign _maxi_read_data_idle = _maxi_read_req_fifo_empty && !_maxi_read_data_busy;
  assign _maxi_read_idle = _maxi_read_req_idle && _maxi_read_data_idle;
  reg _maxi_write_start;
  reg [8-1:0] _maxi_write_op_sel;
  reg [32-1:0] _maxi_write_global_addr;
  reg [33-1:0] _maxi_write_global_size;
  reg [32-1:0] _maxi_write_local_addr;
  reg [32-1:0] _maxi_write_local_stride;
  reg [33-1:0] _maxi_write_local_size;
  reg [32-1:0] _maxi_write_local_blocksize;
  wire _maxi_write_req_fifo_enq;
  wire [137-1:0] _maxi_write_req_fifo_wdata;
  wire _maxi_write_req_fifo_full;
  wire _maxi_write_req_fifo_almost_full;
  wire _maxi_write_req_fifo_deq;
  wire [137-1:0] _maxi_write_req_fifo_rdata;
  wire _maxi_write_req_fifo_empty;
  wire _maxi_write_req_fifo_almost_empty;

  _maxi_write_req_fifo
  inst__maxi_write_req_fifo
  (
    .CLK(CLK),
    .RST(RESETN_inv_buf),
    ._maxi_write_req_fifo_enq(_maxi_write_req_fifo_enq),
    ._maxi_write_req_fifo_wdata(_maxi_write_req_fifo_wdata),
    ._maxi_write_req_fifo_full(_maxi_write_req_fifo_full),
    ._maxi_write_req_fifo_almost_full(_maxi_write_req_fifo_almost_full),
    ._maxi_write_req_fifo_deq(_maxi_write_req_fifo_deq),
    ._maxi_write_req_fifo_rdata(_maxi_write_req_fifo_rdata),
    ._maxi_write_req_fifo_empty(_maxi_write_req_fifo_empty),
    ._maxi_write_req_fifo_almost_empty(_maxi_write_req_fifo_almost_empty)
  );

  reg [4-1:0] count__maxi_write_req_fifo;
  wire [8-1:0] _maxi_write_op_sel_fifo;
  wire [32-1:0] _maxi_write_local_addr_fifo;
  wire [32-1:0] _maxi_write_local_stride_fifo;
  wire [33-1:0] _maxi_write_size_fifo;
  wire [32-1:0] _maxi_write_local_blocksize_fifo;
  wire [8-1:0] unpack_write_req_op_sel_35;
  wire [32-1:0] unpack_write_req_local_addr_36;
  wire [32-1:0] unpack_write_req_local_stride_37;
  wire [33-1:0] unpack_write_req_size_38;
  wire [32-1:0] unpack_write_req_local_blocksize_39;
  assign unpack_write_req_op_sel_35 = _maxi_write_req_fifo_rdata[136:129];
  assign unpack_write_req_local_addr_36 = _maxi_write_req_fifo_rdata[128:97];
  assign unpack_write_req_local_stride_37 = _maxi_write_req_fifo_rdata[96:65];
  assign unpack_write_req_size_38 = _maxi_write_req_fifo_rdata[64:32];
  assign unpack_write_req_local_blocksize_39 = _maxi_write_req_fifo_rdata[31:0];
  assign _maxi_write_op_sel_fifo = unpack_write_req_op_sel_35;
  assign _maxi_write_local_addr_fifo = unpack_write_req_local_addr_36;
  assign _maxi_write_local_stride_fifo = unpack_write_req_local_stride_37;
  assign _maxi_write_size_fifo = unpack_write_req_size_38;
  assign _maxi_write_local_blocksize_fifo = unpack_write_req_local_blocksize_39;
  reg [8-1:0] _maxi_write_op_sel_buf;
  reg [32-1:0] _maxi_write_local_addr_buf;
  reg [32-1:0] _maxi_write_local_stride_buf;
  reg [33-1:0] _maxi_write_size_buf;
  reg [32-1:0] _maxi_write_local_blocksize_buf;
  reg _maxi_write_req_busy;
  reg _maxi_write_data_busy;
  wire _maxi_write_req_idle;
  wire _maxi_write_data_idle;
  wire _maxi_write_idle;
  assign _maxi_write_req_idle = !_maxi_write_start && !_maxi_write_req_busy;
  assign _maxi_write_data_idle = _maxi_write_req_fifo_empty && !_maxi_write_data_busy;
  assign _maxi_write_idle = _maxi_write_req_idle && _maxi_write_data_idle;
  reg [32-1:0] _maxi_global_base_addr;
  assign saxi_bresp = 0;
  assign saxi_rresp = 0;
  reg signed [32-1:0] _saxi_register_0;
  reg signed [32-1:0] _saxi_register_1;
  reg signed [32-1:0] _saxi_register_2;
  reg signed [32-1:0] _saxi_register_3;
  reg signed [32-1:0] _saxi_register_4;
  reg signed [32-1:0] _saxi_register_5;
  reg signed [32-1:0] _saxi_register_6;
  reg signed [32-1:0] _saxi_register_7;
  reg signed [32-1:0] _saxi_register_8;
  reg signed [32-1:0] _saxi_register_9;
  reg signed [32-1:0] _saxi_register_10;
  reg signed [32-1:0] _saxi_register_11;
  reg signed [32-1:0] _saxi_register_12;
  reg signed [32-1:0] _saxi_register_13;
  reg signed [32-1:0] _saxi_register_14;
  reg signed [32-1:0] _saxi_register_15;
  reg signed [32-1:0] _saxi_register_16;
  reg signed [32-1:0] _saxi_register_17;
  reg signed [32-1:0] _saxi_register_18;
  reg signed [32-1:0] _saxi_register_19;
  reg signed [32-1:0] _saxi_register_20;
  reg signed [32-1:0] _saxi_register_21;
  reg signed [32-1:0] _saxi_register_22;
  reg signed [32-1:0] _saxi_register_23;
  reg signed [32-1:0] _saxi_register_24;
  reg signed [32-1:0] _saxi_register_25;
  reg signed [32-1:0] _saxi_register_26;
  reg signed [32-1:0] _saxi_register_27;
  reg signed [32-1:0] _saxi_register_28;
  reg signed [32-1:0] _saxi_register_29;
  reg signed [32-1:0] _saxi_register_30;
  reg signed [32-1:0] _saxi_register_31;
  reg signed [32-1:0] _saxi_register_32;
  reg signed [32-1:0] _saxi_register_33;
  reg signed [32-1:0] _saxi_register_34;
  reg signed [32-1:0] _saxi_register_35;
  reg signed [32-1:0] _saxi_register_36;
  reg _saxi_flag_0;
  reg _saxi_flag_1;
  reg _saxi_flag_2;
  reg _saxi_flag_3;
  reg _saxi_flag_4;
  reg _saxi_flag_5;
  reg _saxi_flag_6;
  reg _saxi_flag_7;
  reg _saxi_flag_8;
  reg _saxi_flag_9;
  reg _saxi_flag_10;
  reg _saxi_flag_11;
  reg _saxi_flag_12;
  reg _saxi_flag_13;
  reg _saxi_flag_14;
  reg _saxi_flag_15;
  reg _saxi_flag_16;
  reg _saxi_flag_17;
  reg _saxi_flag_18;
  reg _saxi_flag_19;
  reg _saxi_flag_20;
  reg _saxi_flag_21;
  reg _saxi_flag_22;
  reg _saxi_flag_23;
  reg _saxi_flag_24;
  reg _saxi_flag_25;
  reg _saxi_flag_26;
  reg _saxi_flag_27;
  reg _saxi_flag_28;
  reg _saxi_flag_29;
  reg _saxi_flag_30;
  reg _saxi_flag_31;
  reg _saxi_flag_32;
  reg _saxi_flag_33;
  reg _saxi_flag_34;
  reg _saxi_flag_35;
  reg _saxi_flag_36;
  reg signed [32-1:0] _saxi_resetval_0;
  reg signed [32-1:0] _saxi_resetval_1;
  reg signed [32-1:0] _saxi_resetval_2;
  reg signed [32-1:0] _saxi_resetval_3;
  reg signed [32-1:0] _saxi_resetval_4;
  reg signed [32-1:0] _saxi_resetval_5;
  reg signed [32-1:0] _saxi_resetval_6;
  reg signed [32-1:0] _saxi_resetval_7;
  reg signed [32-1:0] _saxi_resetval_8;
  reg signed [32-1:0] _saxi_resetval_9;
  reg signed [32-1:0] _saxi_resetval_10;
  reg signed [32-1:0] _saxi_resetval_11;
  reg signed [32-1:0] _saxi_resetval_12;
  reg signed [32-1:0] _saxi_resetval_13;
  reg signed [32-1:0] _saxi_resetval_14;
  reg signed [32-1:0] _saxi_resetval_15;
  reg signed [32-1:0] _saxi_resetval_16;
  reg signed [32-1:0] _saxi_resetval_17;
  reg signed [32-1:0] _saxi_resetval_18;
  reg signed [32-1:0] _saxi_resetval_19;
  reg signed [32-1:0] _saxi_resetval_20;
  reg signed [32-1:0] _saxi_resetval_21;
  reg signed [32-1:0] _saxi_resetval_22;
  reg signed [32-1:0] _saxi_resetval_23;
  reg signed [32-1:0] _saxi_resetval_24;
  reg signed [32-1:0] _saxi_resetval_25;
  reg signed [32-1:0] _saxi_resetval_26;
  reg signed [32-1:0] _saxi_resetval_27;
  reg signed [32-1:0] _saxi_resetval_28;
  reg signed [32-1:0] _saxi_resetval_29;
  reg signed [32-1:0] _saxi_resetval_30;
  reg signed [32-1:0] _saxi_resetval_31;
  reg signed [32-1:0] _saxi_resetval_32;
  reg signed [32-1:0] _saxi_resetval_33;
  reg signed [32-1:0] _saxi_resetval_34;
  reg signed [32-1:0] _saxi_resetval_35;
  reg signed [32-1:0] _saxi_resetval_36;
  localparam _saxi_maskwidth = 6;
  localparam _saxi_mask = { _saxi_maskwidth{ 1'd1 } };
  localparam _saxi_shift = 2;
  reg [32-1:0] _saxi_register_fsm;
  localparam _saxi_register_fsm_init = 0;
  reg [32-1:0] addr_40;
  reg writevalid_41;
  reg readvalid_42;
  reg prev_awvalid_43;
  reg prev_arvalid_44;
  assign saxi_awready = (_saxi_register_fsm == 0) && (!writevalid_41 && !readvalid_42 && !saxi_bvalid && prev_awvalid_43);
  assign saxi_arready = (_saxi_register_fsm == 0) && (!readvalid_42 && !writevalid_41 && prev_arvalid_44 && !prev_awvalid_43);
  reg [_saxi_maskwidth-1:0] axis_maskaddr_45;
  wire signed [32-1:0] axislite_rdata_46;
  assign axislite_rdata_46 = (axis_maskaddr_45 == 0)? _saxi_register_0 : 
                             (axis_maskaddr_45 == 1)? _saxi_register_1 : 
                             (axis_maskaddr_45 == 2)? _saxi_register_2 : 
                             (axis_maskaddr_45 == 3)? _saxi_register_3 : 
                             (axis_maskaddr_45 == 4)? _saxi_register_4 : 
                             (axis_maskaddr_45 == 5)? _saxi_register_5 : 
                             (axis_maskaddr_45 == 6)? _saxi_register_6 : 
                             (axis_maskaddr_45 == 7)? _saxi_register_7 : 
                             (axis_maskaddr_45 == 8)? _saxi_register_8 : 
                             (axis_maskaddr_45 == 9)? _saxi_register_9 : 
                             (axis_maskaddr_45 == 10)? _saxi_register_10 : 
                             (axis_maskaddr_45 == 11)? _saxi_register_11 : 
                             (axis_maskaddr_45 == 12)? _saxi_register_12 : 
                             (axis_maskaddr_45 == 13)? _saxi_register_13 : 
                             (axis_maskaddr_45 == 14)? _saxi_register_14 : 
                             (axis_maskaddr_45 == 15)? _saxi_register_15 : 
                             (axis_maskaddr_45 == 16)? _saxi_register_16 : 
                             (axis_maskaddr_45 == 17)? _saxi_register_17 : 
                             (axis_maskaddr_45 == 18)? _saxi_register_18 : 
                             (axis_maskaddr_45 == 19)? _saxi_register_19 : 
                             (axis_maskaddr_45 == 20)? _saxi_register_20 : 
                             (axis_maskaddr_45 == 21)? _saxi_register_21 : 
                             (axis_maskaddr_45 == 22)? _saxi_register_22 : 
                             (axis_maskaddr_45 == 23)? _saxi_register_23 : 
                             (axis_maskaddr_45 == 24)? _saxi_register_24 : 
                             (axis_maskaddr_45 == 25)? _saxi_register_25 : 
                             (axis_maskaddr_45 == 26)? _saxi_register_26 : 
                             (axis_maskaddr_45 == 27)? _saxi_register_27 : 
                             (axis_maskaddr_45 == 28)? _saxi_register_28 : 
                             (axis_maskaddr_45 == 29)? _saxi_register_29 : 
                             (axis_maskaddr_45 == 30)? _saxi_register_30 : 
                             (axis_maskaddr_45 == 31)? _saxi_register_31 : 
                             (axis_maskaddr_45 == 32)? _saxi_register_32 : 
                             (axis_maskaddr_45 == 33)? _saxi_register_33 : 
                             (axis_maskaddr_45 == 34)? _saxi_register_34 : 
                             (axis_maskaddr_45 == 35)? _saxi_register_35 : 
                             (axis_maskaddr_45 == 36)? _saxi_register_36 : 'hx;
  wire axislite_flag_47;
  assign axislite_flag_47 = (axis_maskaddr_45 == 0)? _saxi_flag_0 : 
                            (axis_maskaddr_45 == 1)? _saxi_flag_1 : 
                            (axis_maskaddr_45 == 2)? _saxi_flag_2 : 
                            (axis_maskaddr_45 == 3)? _saxi_flag_3 : 
                            (axis_maskaddr_45 == 4)? _saxi_flag_4 : 
                            (axis_maskaddr_45 == 5)? _saxi_flag_5 : 
                            (axis_maskaddr_45 == 6)? _saxi_flag_6 : 
                            (axis_maskaddr_45 == 7)? _saxi_flag_7 : 
                            (axis_maskaddr_45 == 8)? _saxi_flag_8 : 
                            (axis_maskaddr_45 == 9)? _saxi_flag_9 : 
                            (axis_maskaddr_45 == 10)? _saxi_flag_10 : 
                            (axis_maskaddr_45 == 11)? _saxi_flag_11 : 
                            (axis_maskaddr_45 == 12)? _saxi_flag_12 : 
                            (axis_maskaddr_45 == 13)? _saxi_flag_13 : 
                            (axis_maskaddr_45 == 14)? _saxi_flag_14 : 
                            (axis_maskaddr_45 == 15)? _saxi_flag_15 : 
                            (axis_maskaddr_45 == 16)? _saxi_flag_16 : 
                            (axis_maskaddr_45 == 17)? _saxi_flag_17 : 
                            (axis_maskaddr_45 == 18)? _saxi_flag_18 : 
                            (axis_maskaddr_45 == 19)? _saxi_flag_19 : 
                            (axis_maskaddr_45 == 20)? _saxi_flag_20 : 
                            (axis_maskaddr_45 == 21)? _saxi_flag_21 : 
                            (axis_maskaddr_45 == 22)? _saxi_flag_22 : 
                            (axis_maskaddr_45 == 23)? _saxi_flag_23 : 
                            (axis_maskaddr_45 == 24)? _saxi_flag_24 : 
                            (axis_maskaddr_45 == 25)? _saxi_flag_25 : 
                            (axis_maskaddr_45 == 26)? _saxi_flag_26 : 
                            (axis_maskaddr_45 == 27)? _saxi_flag_27 : 
                            (axis_maskaddr_45 == 28)? _saxi_flag_28 : 
                            (axis_maskaddr_45 == 29)? _saxi_flag_29 : 
                            (axis_maskaddr_45 == 30)? _saxi_flag_30 : 
                            (axis_maskaddr_45 == 31)? _saxi_flag_31 : 
                            (axis_maskaddr_45 == 32)? _saxi_flag_32 : 
                            (axis_maskaddr_45 == 33)? _saxi_flag_33 : 
                            (axis_maskaddr_45 == 34)? _saxi_flag_34 : 
                            (axis_maskaddr_45 == 35)? _saxi_flag_35 : 
                            (axis_maskaddr_45 == 36)? _saxi_flag_36 : 'hx;
  wire signed [32-1:0] axislite_resetval_48;
  assign axislite_resetval_48 = (axis_maskaddr_45 == 0)? _saxi_resetval_0 : 
                                (axis_maskaddr_45 == 1)? _saxi_resetval_1 : 
                                (axis_maskaddr_45 == 2)? _saxi_resetval_2 : 
                                (axis_maskaddr_45 == 3)? _saxi_resetval_3 : 
                                (axis_maskaddr_45 == 4)? _saxi_resetval_4 : 
                                (axis_maskaddr_45 == 5)? _saxi_resetval_5 : 
                                (axis_maskaddr_45 == 6)? _saxi_resetval_6 : 
                                (axis_maskaddr_45 == 7)? _saxi_resetval_7 : 
                                (axis_maskaddr_45 == 8)? _saxi_resetval_8 : 
                                (axis_maskaddr_45 == 9)? _saxi_resetval_9 : 
                                (axis_maskaddr_45 == 10)? _saxi_resetval_10 : 
                                (axis_maskaddr_45 == 11)? _saxi_resetval_11 : 
                                (axis_maskaddr_45 == 12)? _saxi_resetval_12 : 
                                (axis_maskaddr_45 == 13)? _saxi_resetval_13 : 
                                (axis_maskaddr_45 == 14)? _saxi_resetval_14 : 
                                (axis_maskaddr_45 == 15)? _saxi_resetval_15 : 
                                (axis_maskaddr_45 == 16)? _saxi_resetval_16 : 
                                (axis_maskaddr_45 == 17)? _saxi_resetval_17 : 
                                (axis_maskaddr_45 == 18)? _saxi_resetval_18 : 
                                (axis_maskaddr_45 == 19)? _saxi_resetval_19 : 
                                (axis_maskaddr_45 == 20)? _saxi_resetval_20 : 
                                (axis_maskaddr_45 == 21)? _saxi_resetval_21 : 
                                (axis_maskaddr_45 == 22)? _saxi_resetval_22 : 
                                (axis_maskaddr_45 == 23)? _saxi_resetval_23 : 
                                (axis_maskaddr_45 == 24)? _saxi_resetval_24 : 
                                (axis_maskaddr_45 == 25)? _saxi_resetval_25 : 
                                (axis_maskaddr_45 == 26)? _saxi_resetval_26 : 
                                (axis_maskaddr_45 == 27)? _saxi_resetval_27 : 
                                (axis_maskaddr_45 == 28)? _saxi_resetval_28 : 
                                (axis_maskaddr_45 == 29)? _saxi_resetval_29 : 
                                (axis_maskaddr_45 == 30)? _saxi_resetval_30 : 
                                (axis_maskaddr_45 == 31)? _saxi_resetval_31 : 
                                (axis_maskaddr_45 == 32)? _saxi_resetval_32 : 
                                (axis_maskaddr_45 == 33)? _saxi_resetval_33 : 
                                (axis_maskaddr_45 == 34)? _saxi_resetval_34 : 
                                (axis_maskaddr_45 == 35)? _saxi_resetval_35 : 
                                (axis_maskaddr_45 == 36)? _saxi_resetval_36 : 'hx;
  reg _saxi_rdata_cond_0_1;
  assign saxi_wready = _saxi_register_fsm == 3;
  wire maxi_idle;
  assign maxi_idle = _maxi_write_idle & _maxi_read_idle;
  wire sw_rst_logic;
  assign sw_rst_logic = maxi_idle & _saxi_register_6;
  wire rst_logic;
  assign rst_logic = RESETN_inv_buf | sw_rst_logic;
  reg RST;
  reg _rst_logic_1;
  reg _rst_logic_2;
  wire signed [32-1:0] irq_49;
  assign irq_49 = _saxi_register_9 & _saxi_register_10;
  wire irq_busy;
  assign irq_busy = _saxi_register_5[0];
  reg irq_busy_edge_50;
  wire irq_busy_edge_51;
  assign irq_busy_edge_51 = irq_busy_edge_50 & !irq_busy;
  wire irq_extern;
  assign irq_extern = |_saxi_register_7;
  reg irq_extern_edge_52;
  wire irq_extern_edge_53;
  assign irq_extern_edge_53 = !irq_extern_edge_52 & irq_extern;
  wire [15-1:0] ram_w32_l32768_id0_0_addr;
  wire [32-1:0] ram_w32_l32768_id0_0_rdata;
  wire [32-1:0] ram_w32_l32768_id0_0_wdata;
  wire ram_w32_l32768_id0_0_wenable;
  wire ram_w32_l32768_id0_0_enable;
  wire [15-1:0] ram_w32_l32768_id0_1_addr;
  wire [32-1:0] ram_w32_l32768_id0_1_rdata;
  wire [32-1:0] ram_w32_l32768_id0_1_wdata;
  wire ram_w32_l32768_id0_1_wenable;
  wire ram_w32_l32768_id0_1_enable;
  assign ram_w32_l32768_id0_0_wdata = 'hx;
  assign ram_w32_l32768_id0_0_wenable = 0;

  ram_w32_l32768_id0
  inst_ram_w32_l32768_id0
  (
    .CLK(CLK),
    .ram_w32_l32768_id0_0_addr(ram_w32_l32768_id0_0_addr),
    .ram_w32_l32768_id0_0_rdata(ram_w32_l32768_id0_0_rdata),
    .ram_w32_l32768_id0_0_wdata(ram_w32_l32768_id0_0_wdata),
    .ram_w32_l32768_id0_0_wenable(ram_w32_l32768_id0_0_wenable),
    .ram_w32_l32768_id0_0_enable(ram_w32_l32768_id0_0_enable),
    .ram_w32_l32768_id0_1_addr(ram_w32_l32768_id0_1_addr),
    .ram_w32_l32768_id0_1_rdata(ram_w32_l32768_id0_1_rdata),
    .ram_w32_l32768_id0_1_wdata(ram_w32_l32768_id0_1_wdata),
    .ram_w32_l32768_id0_1_wenable(ram_w32_l32768_id0_1_wenable),
    .ram_w32_l32768_id0_1_enable(ram_w32_l32768_id0_1_enable)
  );

  wire [14-1:0] ram_w32_l16384_id0_0_addr;
  wire [32-1:0] ram_w32_l16384_id0_0_rdata;
  wire [32-1:0] ram_w32_l16384_id0_0_wdata;
  wire ram_w32_l16384_id0_0_wenable;
  wire ram_w32_l16384_id0_0_enable;
  wire [14-1:0] ram_w32_l16384_id0_1_addr;
  wire [32-1:0] ram_w32_l16384_id0_1_rdata;
  wire [32-1:0] ram_w32_l16384_id0_1_wdata;
  wire ram_w32_l16384_id0_1_wenable;
  wire ram_w32_l16384_id0_1_enable;
  assign ram_w32_l16384_id0_1_wdata = 'hx;
  assign ram_w32_l16384_id0_1_wenable = 0;

  ram_w32_l16384_id0
  inst_ram_w32_l16384_id0
  (
    .CLK(CLK),
    .ram_w32_l16384_id0_0_addr(ram_w32_l16384_id0_0_addr),
    .ram_w32_l16384_id0_0_rdata(ram_w32_l16384_id0_0_rdata),
    .ram_w32_l16384_id0_0_wdata(ram_w32_l16384_id0_0_wdata),
    .ram_w32_l16384_id0_0_wenable(ram_w32_l16384_id0_0_wenable),
    .ram_w32_l16384_id0_0_enable(ram_w32_l16384_id0_0_enable),
    .ram_w32_l16384_id0_1_addr(ram_w32_l16384_id0_1_addr),
    .ram_w32_l16384_id0_1_rdata(ram_w32_l16384_id0_1_rdata),
    .ram_w32_l16384_id0_1_wdata(ram_w32_l16384_id0_1_wdata),
    .ram_w32_l16384_id0_1_wenable(ram_w32_l16384_id0_1_wenable),
    .ram_w32_l16384_id0_1_enable(ram_w32_l16384_id0_1_enable)
  );

  wire [13-1:0] ram_w32_l8192_id0_0_addr;
  wire [32-1:0] ram_w32_l8192_id0_0_rdata;
  wire [32-1:0] ram_w32_l8192_id0_0_wdata;
  wire ram_w32_l8192_id0_0_wenable;
  wire ram_w32_l8192_id0_0_enable;
  wire [13-1:0] ram_w32_l8192_id0_1_addr;
  wire [32-1:0] ram_w32_l8192_id0_1_rdata;
  wire [32-1:0] ram_w32_l8192_id0_1_wdata;
  wire ram_w32_l8192_id0_1_wenable;
  wire ram_w32_l8192_id0_1_enable;

  ram_w32_l8192_id0
  inst_ram_w32_l8192_id0
  (
    .CLK(CLK),
    .ram_w32_l8192_id0_0_addr(ram_w32_l8192_id0_0_addr),
    .ram_w32_l8192_id0_0_rdata(ram_w32_l8192_id0_0_rdata),
    .ram_w32_l8192_id0_0_wdata(ram_w32_l8192_id0_0_wdata),
    .ram_w32_l8192_id0_0_wenable(ram_w32_l8192_id0_0_wenable),
    .ram_w32_l8192_id0_0_enable(ram_w32_l8192_id0_0_enable),
    .ram_w32_l8192_id0_1_addr(ram_w32_l8192_id0_1_addr),
    .ram_w32_l8192_id0_1_rdata(ram_w32_l8192_id0_1_rdata),
    .ram_w32_l8192_id0_1_wdata(ram_w32_l8192_id0_1_wdata),
    .ram_w32_l8192_id0_1_wenable(ram_w32_l8192_id0_1_wenable),
    .ram_w32_l8192_id0_1_enable(ram_w32_l8192_id0_1_enable)
  );

  wire [13-1:0] ram_w32_l8192_id1_0_addr;
  wire [32-1:0] ram_w32_l8192_id1_0_rdata;
  wire [32-1:0] ram_w32_l8192_id1_0_wdata;
  wire ram_w32_l8192_id1_0_wenable;
  wire ram_w32_l8192_id1_0_enable;
  wire [13-1:0] ram_w32_l8192_id1_1_addr;
  wire [32-1:0] ram_w32_l8192_id1_1_rdata;
  wire [32-1:0] ram_w32_l8192_id1_1_wdata;
  wire ram_w32_l8192_id1_1_wenable;
  wire ram_w32_l8192_id1_1_enable;
  assign ram_w32_l8192_id1_0_wdata = 'hx;
  assign ram_w32_l8192_id1_0_wenable = 0;

  ram_w32_l8192_id1
  inst_ram_w32_l8192_id1
  (
    .CLK(CLK),
    .ram_w32_l8192_id1_0_addr(ram_w32_l8192_id1_0_addr),
    .ram_w32_l8192_id1_0_rdata(ram_w32_l8192_id1_0_rdata),
    .ram_w32_l8192_id1_0_wdata(ram_w32_l8192_id1_0_wdata),
    .ram_w32_l8192_id1_0_wenable(ram_w32_l8192_id1_0_wenable),
    .ram_w32_l8192_id1_0_enable(ram_w32_l8192_id1_0_enable),
    .ram_w32_l8192_id1_1_addr(ram_w32_l8192_id1_1_addr),
    .ram_w32_l8192_id1_1_rdata(ram_w32_l8192_id1_1_rdata),
    .ram_w32_l8192_id1_1_wdata(ram_w32_l8192_id1_1_wdata),
    .ram_w32_l8192_id1_1_wenable(ram_w32_l8192_id1_1_wenable),
    .ram_w32_l8192_id1_1_enable(ram_w32_l8192_id1_1_enable)
  );

  wire [13-1:0] ram_w32_l8192_id2_0_addr;
  wire [32-1:0] ram_w32_l8192_id2_0_rdata;
  wire [32-1:0] ram_w32_l8192_id2_0_wdata;
  wire ram_w32_l8192_id2_0_wenable;
  wire ram_w32_l8192_id2_0_enable;
  wire [13-1:0] ram_w32_l8192_id2_1_addr;
  wire [32-1:0] ram_w32_l8192_id2_1_rdata;
  wire [32-1:0] ram_w32_l8192_id2_1_wdata;
  wire ram_w32_l8192_id2_1_wenable;
  wire ram_w32_l8192_id2_1_enable;
  assign ram_w32_l8192_id2_0_wdata = 'hx;
  assign ram_w32_l8192_id2_0_wenable = 0;

  ram_w32_l8192_id2
  inst_ram_w32_l8192_id2
  (
    .CLK(CLK),
    .ram_w32_l8192_id2_0_addr(ram_w32_l8192_id2_0_addr),
    .ram_w32_l8192_id2_0_rdata(ram_w32_l8192_id2_0_rdata),
    .ram_w32_l8192_id2_0_wdata(ram_w32_l8192_id2_0_wdata),
    .ram_w32_l8192_id2_0_wenable(ram_w32_l8192_id2_0_wenable),
    .ram_w32_l8192_id2_0_enable(ram_w32_l8192_id2_0_enable),
    .ram_w32_l8192_id2_1_addr(ram_w32_l8192_id2_1_addr),
    .ram_w32_l8192_id2_1_rdata(ram_w32_l8192_id2_1_rdata),
    .ram_w32_l8192_id2_1_wdata(ram_w32_l8192_id2_1_wdata),
    .ram_w32_l8192_id2_1_wenable(ram_w32_l8192_id2_1_wenable),
    .ram_w32_l8192_id2_1_enable(ram_w32_l8192_id2_1_enable)
  );

  wire [13-1:0] ram_w32_l8192_id3_0_addr;
  wire [32-1:0] ram_w32_l8192_id3_0_rdata;
  wire [32-1:0] ram_w32_l8192_id3_0_wdata;
  wire ram_w32_l8192_id3_0_wenable;
  wire ram_w32_l8192_id3_0_enable;
  wire [13-1:0] ram_w32_l8192_id3_1_addr;
  wire [32-1:0] ram_w32_l8192_id3_1_rdata;
  wire [32-1:0] ram_w32_l8192_id3_1_wdata;
  wire ram_w32_l8192_id3_1_wenable;
  wire ram_w32_l8192_id3_1_enable;
  assign ram_w32_l8192_id3_0_wdata = 'hx;
  assign ram_w32_l8192_id3_0_wenable = 0;

  ram_w32_l8192_id3
  inst_ram_w32_l8192_id3
  (
    .CLK(CLK),
    .ram_w32_l8192_id3_0_addr(ram_w32_l8192_id3_0_addr),
    .ram_w32_l8192_id3_0_rdata(ram_w32_l8192_id3_0_rdata),
    .ram_w32_l8192_id3_0_wdata(ram_w32_l8192_id3_0_wdata),
    .ram_w32_l8192_id3_0_wenable(ram_w32_l8192_id3_0_wenable),
    .ram_w32_l8192_id3_0_enable(ram_w32_l8192_id3_0_enable),
    .ram_w32_l8192_id3_1_addr(ram_w32_l8192_id3_1_addr),
    .ram_w32_l8192_id3_1_rdata(ram_w32_l8192_id3_1_rdata),
    .ram_w32_l8192_id3_1_wdata(ram_w32_l8192_id3_1_wdata),
    .ram_w32_l8192_id3_1_wenable(ram_w32_l8192_id3_1_wenable),
    .ram_w32_l8192_id3_1_enable(ram_w32_l8192_id3_1_enable)
  );

  wire [12-1:0] ram_w32_l4096_id0_0_addr;
  wire [32-1:0] ram_w32_l4096_id0_0_rdata;
  wire [32-1:0] ram_w32_l4096_id0_0_wdata;
  wire ram_w32_l4096_id0_0_wenable;
  wire ram_w32_l4096_id0_0_enable;
  wire [12-1:0] ram_w32_l4096_id0_1_addr;
  wire [32-1:0] ram_w32_l4096_id0_1_rdata;
  wire [32-1:0] ram_w32_l4096_id0_1_wdata;
  wire ram_w32_l4096_id0_1_wenable;
  wire ram_w32_l4096_id0_1_enable;
  assign ram_w32_l4096_id0_0_wdata = 'hx;
  assign ram_w32_l4096_id0_0_wenable = 0;

  ram_w32_l4096_id0
  inst_ram_w32_l4096_id0
  (
    .CLK(CLK),
    .ram_w32_l4096_id0_0_addr(ram_w32_l4096_id0_0_addr),
    .ram_w32_l4096_id0_0_rdata(ram_w32_l4096_id0_0_rdata),
    .ram_w32_l4096_id0_0_wdata(ram_w32_l4096_id0_0_wdata),
    .ram_w32_l4096_id0_0_wenable(ram_w32_l4096_id0_0_wenable),
    .ram_w32_l4096_id0_0_enable(ram_w32_l4096_id0_0_enable),
    .ram_w32_l4096_id0_1_addr(ram_w32_l4096_id0_1_addr),
    .ram_w32_l4096_id0_1_rdata(ram_w32_l4096_id0_1_rdata),
    .ram_w32_l4096_id0_1_wdata(ram_w32_l4096_id0_1_wdata),
    .ram_w32_l4096_id0_1_wenable(ram_w32_l4096_id0_1_wenable),
    .ram_w32_l4096_id0_1_enable(ram_w32_l4096_id0_1_enable)
  );

  wire [12-1:0] ram_w32_l4096_id1_0_addr;
  wire [32-1:0] ram_w32_l4096_id1_0_rdata;
  wire [32-1:0] ram_w32_l4096_id1_0_wdata;
  wire ram_w32_l4096_id1_0_wenable;
  wire ram_w32_l4096_id1_0_enable;
  wire [12-1:0] ram_w32_l4096_id1_1_addr;
  wire [32-1:0] ram_w32_l4096_id1_1_rdata;
  wire [32-1:0] ram_w32_l4096_id1_1_wdata;
  wire ram_w32_l4096_id1_1_wenable;
  wire ram_w32_l4096_id1_1_enable;
  assign ram_w32_l4096_id1_0_wdata = 'hx;
  assign ram_w32_l4096_id1_0_wenable = 0;

  ram_w32_l4096_id1
  inst_ram_w32_l4096_id1
  (
    .CLK(CLK),
    .ram_w32_l4096_id1_0_addr(ram_w32_l4096_id1_0_addr),
    .ram_w32_l4096_id1_0_rdata(ram_w32_l4096_id1_0_rdata),
    .ram_w32_l4096_id1_0_wdata(ram_w32_l4096_id1_0_wdata),
    .ram_w32_l4096_id1_0_wenable(ram_w32_l4096_id1_0_wenable),
    .ram_w32_l4096_id1_0_enable(ram_w32_l4096_id1_0_enable),
    .ram_w32_l4096_id1_1_addr(ram_w32_l4096_id1_1_addr),
    .ram_w32_l4096_id1_1_rdata(ram_w32_l4096_id1_1_rdata),
    .ram_w32_l4096_id1_1_wdata(ram_w32_l4096_id1_1_wdata),
    .ram_w32_l4096_id1_1_wenable(ram_w32_l4096_id1_1_wenable),
    .ram_w32_l4096_id1_1_enable(ram_w32_l4096_id1_1_enable)
  );

  wire [12-1:0] ram_w32_l4096_id2_0_addr;
  wire [32-1:0] ram_w32_l4096_id2_0_rdata;
  wire [32-1:0] ram_w32_l4096_id2_0_wdata;
  wire ram_w32_l4096_id2_0_wenable;
  wire ram_w32_l4096_id2_0_enable;
  wire [12-1:0] ram_w32_l4096_id2_1_addr;
  wire [32-1:0] ram_w32_l4096_id2_1_rdata;
  wire [32-1:0] ram_w32_l4096_id2_1_wdata;
  wire ram_w32_l4096_id2_1_wenable;
  wire ram_w32_l4096_id2_1_enable;
  assign ram_w32_l4096_id2_0_wdata = 'hx;
  assign ram_w32_l4096_id2_0_wenable = 0;

  ram_w32_l4096_id2
  inst_ram_w32_l4096_id2
  (
    .CLK(CLK),
    .ram_w32_l4096_id2_0_addr(ram_w32_l4096_id2_0_addr),
    .ram_w32_l4096_id2_0_rdata(ram_w32_l4096_id2_0_rdata),
    .ram_w32_l4096_id2_0_wdata(ram_w32_l4096_id2_0_wdata),
    .ram_w32_l4096_id2_0_wenable(ram_w32_l4096_id2_0_wenable),
    .ram_w32_l4096_id2_0_enable(ram_w32_l4096_id2_0_enable),
    .ram_w32_l4096_id2_1_addr(ram_w32_l4096_id2_1_addr),
    .ram_w32_l4096_id2_1_rdata(ram_w32_l4096_id2_1_rdata),
    .ram_w32_l4096_id2_1_wdata(ram_w32_l4096_id2_1_wdata),
    .ram_w32_l4096_id2_1_wenable(ram_w32_l4096_id2_1_wenable),
    .ram_w32_l4096_id2_1_enable(ram_w32_l4096_id2_1_enable)
  );

  wire [12-1:0] ram_w32_l4096_id3_0_addr;
  wire [32-1:0] ram_w32_l4096_id3_0_rdata;
  wire [32-1:0] ram_w32_l4096_id3_0_wdata;
  wire ram_w32_l4096_id3_0_wenable;
  wire ram_w32_l4096_id3_0_enable;
  wire [12-1:0] ram_w32_l4096_id3_1_addr;
  wire [32-1:0] ram_w32_l4096_id3_1_rdata;
  wire [32-1:0] ram_w32_l4096_id3_1_wdata;
  wire ram_w32_l4096_id3_1_wenable;
  wire ram_w32_l4096_id3_1_enable;
  assign ram_w32_l4096_id3_0_wdata = 'hx;
  assign ram_w32_l4096_id3_0_wenable = 0;

  ram_w32_l4096_id3
  inst_ram_w32_l4096_id3
  (
    .CLK(CLK),
    .ram_w32_l4096_id3_0_addr(ram_w32_l4096_id3_0_addr),
    .ram_w32_l4096_id3_0_rdata(ram_w32_l4096_id3_0_rdata),
    .ram_w32_l4096_id3_0_wdata(ram_w32_l4096_id3_0_wdata),
    .ram_w32_l4096_id3_0_wenable(ram_w32_l4096_id3_0_wenable),
    .ram_w32_l4096_id3_0_enable(ram_w32_l4096_id3_0_enable),
    .ram_w32_l4096_id3_1_addr(ram_w32_l4096_id3_1_addr),
    .ram_w32_l4096_id3_1_rdata(ram_w32_l4096_id3_1_rdata),
    .ram_w32_l4096_id3_1_wdata(ram_w32_l4096_id3_1_wdata),
    .ram_w32_l4096_id3_1_wenable(ram_w32_l4096_id3_1_wenable),
    .ram_w32_l4096_id3_1_enable(ram_w32_l4096_id3_1_enable)
  );

  wire [12-1:0] ram_w32_l4096_id4_0_addr;
  wire [32-1:0] ram_w32_l4096_id4_0_rdata;
  wire [32-1:0] ram_w32_l4096_id4_0_wdata;
  wire ram_w32_l4096_id4_0_wenable;
  wire ram_w32_l4096_id4_0_enable;
  wire [12-1:0] ram_w32_l4096_id4_1_addr;
  wire [32-1:0] ram_w32_l4096_id4_1_rdata;
  wire [32-1:0] ram_w32_l4096_id4_1_wdata;
  wire ram_w32_l4096_id4_1_wenable;
  wire ram_w32_l4096_id4_1_enable;
  assign ram_w32_l4096_id4_0_wdata = 'hx;
  assign ram_w32_l4096_id4_0_wenable = 0;

  ram_w32_l4096_id4
  inst_ram_w32_l4096_id4
  (
    .CLK(CLK),
    .ram_w32_l4096_id4_0_addr(ram_w32_l4096_id4_0_addr),
    .ram_w32_l4096_id4_0_rdata(ram_w32_l4096_id4_0_rdata),
    .ram_w32_l4096_id4_0_wdata(ram_w32_l4096_id4_0_wdata),
    .ram_w32_l4096_id4_0_wenable(ram_w32_l4096_id4_0_wenable),
    .ram_w32_l4096_id4_0_enable(ram_w32_l4096_id4_0_enable),
    .ram_w32_l4096_id4_1_addr(ram_w32_l4096_id4_1_addr),
    .ram_w32_l4096_id4_1_rdata(ram_w32_l4096_id4_1_rdata),
    .ram_w32_l4096_id4_1_wdata(ram_w32_l4096_id4_1_wdata),
    .ram_w32_l4096_id4_1_wenable(ram_w32_l4096_id4_1_wenable),
    .ram_w32_l4096_id4_1_enable(ram_w32_l4096_id4_1_enable)
  );

  wire [12-1:0] ram_w32_l4096_id5_0_addr;
  wire [32-1:0] ram_w32_l4096_id5_0_rdata;
  wire [32-1:0] ram_w32_l4096_id5_0_wdata;
  wire ram_w32_l4096_id5_0_wenable;
  wire ram_w32_l4096_id5_0_enable;
  wire [12-1:0] ram_w32_l4096_id5_1_addr;
  wire [32-1:0] ram_w32_l4096_id5_1_rdata;
  wire [32-1:0] ram_w32_l4096_id5_1_wdata;
  wire ram_w32_l4096_id5_1_wenable;
  wire ram_w32_l4096_id5_1_enable;
  assign ram_w32_l4096_id5_0_wdata = 'hx;
  assign ram_w32_l4096_id5_0_wenable = 0;

  ram_w32_l4096_id5
  inst_ram_w32_l4096_id5
  (
    .CLK(CLK),
    .ram_w32_l4096_id5_0_addr(ram_w32_l4096_id5_0_addr),
    .ram_w32_l4096_id5_0_rdata(ram_w32_l4096_id5_0_rdata),
    .ram_w32_l4096_id5_0_wdata(ram_w32_l4096_id5_0_wdata),
    .ram_w32_l4096_id5_0_wenable(ram_w32_l4096_id5_0_wenable),
    .ram_w32_l4096_id5_0_enable(ram_w32_l4096_id5_0_enable),
    .ram_w32_l4096_id5_1_addr(ram_w32_l4096_id5_1_addr),
    .ram_w32_l4096_id5_1_rdata(ram_w32_l4096_id5_1_rdata),
    .ram_w32_l4096_id5_1_wdata(ram_w32_l4096_id5_1_wdata),
    .ram_w32_l4096_id5_1_wenable(ram_w32_l4096_id5_1_wenable),
    .ram_w32_l4096_id5_1_enable(ram_w32_l4096_id5_1_enable)
  );

  wire [12-1:0] ram_w32_l4096_id6_0_addr;
  wire [32-1:0] ram_w32_l4096_id6_0_rdata;
  wire [32-1:0] ram_w32_l4096_id6_0_wdata;
  wire ram_w32_l4096_id6_0_wenable;
  wire ram_w32_l4096_id6_0_enable;
  wire [12-1:0] ram_w32_l4096_id6_1_addr;
  wire [32-1:0] ram_w32_l4096_id6_1_rdata;
  wire [32-1:0] ram_w32_l4096_id6_1_wdata;
  wire ram_w32_l4096_id6_1_wenable;
  wire ram_w32_l4096_id6_1_enable;
  assign ram_w32_l4096_id6_0_wdata = 'hx;
  assign ram_w32_l4096_id6_0_wenable = 0;

  ram_w32_l4096_id6
  inst_ram_w32_l4096_id6
  (
    .CLK(CLK),
    .ram_w32_l4096_id6_0_addr(ram_w32_l4096_id6_0_addr),
    .ram_w32_l4096_id6_0_rdata(ram_w32_l4096_id6_0_rdata),
    .ram_w32_l4096_id6_0_wdata(ram_w32_l4096_id6_0_wdata),
    .ram_w32_l4096_id6_0_wenable(ram_w32_l4096_id6_0_wenable),
    .ram_w32_l4096_id6_0_enable(ram_w32_l4096_id6_0_enable),
    .ram_w32_l4096_id6_1_addr(ram_w32_l4096_id6_1_addr),
    .ram_w32_l4096_id6_1_rdata(ram_w32_l4096_id6_1_rdata),
    .ram_w32_l4096_id6_1_wdata(ram_w32_l4096_id6_1_wdata),
    .ram_w32_l4096_id6_1_wenable(ram_w32_l4096_id6_1_wenable),
    .ram_w32_l4096_id6_1_enable(ram_w32_l4096_id6_1_enable)
  );

  wire [12-1:0] ram_w32_l4096_id7_0_addr;
  wire [32-1:0] ram_w32_l4096_id7_0_rdata;
  wire [32-1:0] ram_w32_l4096_id7_0_wdata;
  wire ram_w32_l4096_id7_0_wenable;
  wire ram_w32_l4096_id7_0_enable;
  wire [12-1:0] ram_w32_l4096_id7_1_addr;
  wire [32-1:0] ram_w32_l4096_id7_1_rdata;
  wire [32-1:0] ram_w32_l4096_id7_1_wdata;
  wire ram_w32_l4096_id7_1_wenable;
  wire ram_w32_l4096_id7_1_enable;
  assign ram_w32_l4096_id7_0_wdata = 'hx;
  assign ram_w32_l4096_id7_0_wenable = 0;

  ram_w32_l4096_id7
  inst_ram_w32_l4096_id7
  (
    .CLK(CLK),
    .ram_w32_l4096_id7_0_addr(ram_w32_l4096_id7_0_addr),
    .ram_w32_l4096_id7_0_rdata(ram_w32_l4096_id7_0_rdata),
    .ram_w32_l4096_id7_0_wdata(ram_w32_l4096_id7_0_wdata),
    .ram_w32_l4096_id7_0_wenable(ram_w32_l4096_id7_0_wenable),
    .ram_w32_l4096_id7_0_enable(ram_w32_l4096_id7_0_enable),
    .ram_w32_l4096_id7_1_addr(ram_w32_l4096_id7_1_addr),
    .ram_w32_l4096_id7_1_rdata(ram_w32_l4096_id7_1_rdata),
    .ram_w32_l4096_id7_1_wdata(ram_w32_l4096_id7_1_wdata),
    .ram_w32_l4096_id7_1_wenable(ram_w32_l4096_id7_1_wenable),
    .ram_w32_l4096_id7_1_enable(ram_w32_l4096_id7_1_enable)
  );

  wire [12-1:0] ram_w32_l4096_id8_0_addr;
  wire [32-1:0] ram_w32_l4096_id8_0_rdata;
  wire [32-1:0] ram_w32_l4096_id8_0_wdata;
  wire ram_w32_l4096_id8_0_wenable;
  wire ram_w32_l4096_id8_0_enable;
  wire [12-1:0] ram_w32_l4096_id8_1_addr;
  wire [32-1:0] ram_w32_l4096_id8_1_rdata;
  wire [32-1:0] ram_w32_l4096_id8_1_wdata;
  wire ram_w32_l4096_id8_1_wenable;
  wire ram_w32_l4096_id8_1_enable;
  assign ram_w32_l4096_id8_0_wdata = 'hx;
  assign ram_w32_l4096_id8_0_wenable = 0;

  ram_w32_l4096_id8
  inst_ram_w32_l4096_id8
  (
    .CLK(CLK),
    .ram_w32_l4096_id8_0_addr(ram_w32_l4096_id8_0_addr),
    .ram_w32_l4096_id8_0_rdata(ram_w32_l4096_id8_0_rdata),
    .ram_w32_l4096_id8_0_wdata(ram_w32_l4096_id8_0_wdata),
    .ram_w32_l4096_id8_0_wenable(ram_w32_l4096_id8_0_wenable),
    .ram_w32_l4096_id8_0_enable(ram_w32_l4096_id8_0_enable),
    .ram_w32_l4096_id8_1_addr(ram_w32_l4096_id8_1_addr),
    .ram_w32_l4096_id8_1_rdata(ram_w32_l4096_id8_1_rdata),
    .ram_w32_l4096_id8_1_wdata(ram_w32_l4096_id8_1_wdata),
    .ram_w32_l4096_id8_1_wenable(ram_w32_l4096_id8_1_wenable),
    .ram_w32_l4096_id8_1_enable(ram_w32_l4096_id8_1_enable)
  );

  wire [10-1:0] ram_w32_l1024_id0_0_addr;
  wire [32-1:0] ram_w32_l1024_id0_0_rdata;
  wire [32-1:0] ram_w32_l1024_id0_0_wdata;
  wire ram_w32_l1024_id0_0_wenable;
  wire ram_w32_l1024_id0_0_enable;
  wire [10-1:0] ram_w32_l1024_id0_1_addr;
  wire [32-1:0] ram_w32_l1024_id0_1_rdata;
  wire [32-1:0] ram_w32_l1024_id0_1_wdata;
  wire ram_w32_l1024_id0_1_wenable;
  wire ram_w32_l1024_id0_1_enable;
  assign ram_w32_l1024_id0_0_wdata = 'hx;
  assign ram_w32_l1024_id0_0_wenable = 0;

  ram_w32_l1024_id0
  inst_ram_w32_l1024_id0
  (
    .CLK(CLK),
    .ram_w32_l1024_id0_0_addr(ram_w32_l1024_id0_0_addr),
    .ram_w32_l1024_id0_0_rdata(ram_w32_l1024_id0_0_rdata),
    .ram_w32_l1024_id0_0_wdata(ram_w32_l1024_id0_0_wdata),
    .ram_w32_l1024_id0_0_wenable(ram_w32_l1024_id0_0_wenable),
    .ram_w32_l1024_id0_0_enable(ram_w32_l1024_id0_0_enable),
    .ram_w32_l1024_id0_1_addr(ram_w32_l1024_id0_1_addr),
    .ram_w32_l1024_id0_1_rdata(ram_w32_l1024_id0_1_rdata),
    .ram_w32_l1024_id0_1_wdata(ram_w32_l1024_id0_1_wdata),
    .ram_w32_l1024_id0_1_wenable(ram_w32_l1024_id0_1_wenable),
    .ram_w32_l1024_id0_1_enable(ram_w32_l1024_id0_1_enable)
  );

  wire [10-1:0] ram_w32_l1024_id1_0_addr;
  wire [32-1:0] ram_w32_l1024_id1_0_rdata;
  wire [32-1:0] ram_w32_l1024_id1_0_wdata;
  wire ram_w32_l1024_id1_0_wenable;
  wire ram_w32_l1024_id1_0_enable;
  wire [10-1:0] ram_w32_l1024_id1_1_addr;
  wire [32-1:0] ram_w32_l1024_id1_1_rdata;
  wire [32-1:0] ram_w32_l1024_id1_1_wdata;
  wire ram_w32_l1024_id1_1_wenable;
  wire ram_w32_l1024_id1_1_enable;
  assign ram_w32_l1024_id1_1_wdata = 'hx;
  assign ram_w32_l1024_id1_1_wenable = 0;

  ram_w32_l1024_id1
  inst_ram_w32_l1024_id1
  (
    .CLK(CLK),
    .ram_w32_l1024_id1_0_addr(ram_w32_l1024_id1_0_addr),
    .ram_w32_l1024_id1_0_rdata(ram_w32_l1024_id1_0_rdata),
    .ram_w32_l1024_id1_0_wdata(ram_w32_l1024_id1_0_wdata),
    .ram_w32_l1024_id1_0_wenable(ram_w32_l1024_id1_0_wenable),
    .ram_w32_l1024_id1_0_enable(ram_w32_l1024_id1_0_enable),
    .ram_w32_l1024_id1_1_addr(ram_w32_l1024_id1_1_addr),
    .ram_w32_l1024_id1_1_rdata(ram_w32_l1024_id1_1_rdata),
    .ram_w32_l1024_id1_1_wdata(ram_w32_l1024_id1_1_wdata),
    .ram_w32_l1024_id1_1_wenable(ram_w32_l1024_id1_1_wenable),
    .ram_w32_l1024_id1_1_enable(ram_w32_l1024_id1_1_enable)
  );

  wire [10-1:0] ram_w32_l1024_id2_0_addr;
  wire [32-1:0] ram_w32_l1024_id2_0_rdata;
  wire [32-1:0] ram_w32_l1024_id2_0_wdata;
  wire ram_w32_l1024_id2_0_wenable;
  wire ram_w32_l1024_id2_0_enable;
  wire [10-1:0] ram_w32_l1024_id2_1_addr;
  wire [32-1:0] ram_w32_l1024_id2_1_rdata;
  wire [32-1:0] ram_w32_l1024_id2_1_wdata;
  wire ram_w32_l1024_id2_1_wenable;
  wire ram_w32_l1024_id2_1_enable;
  assign ram_w32_l1024_id2_0_wdata = 'hx;
  assign ram_w32_l1024_id2_0_wenable = 0;

  ram_w32_l1024_id2
  inst_ram_w32_l1024_id2
  (
    .CLK(CLK),
    .ram_w32_l1024_id2_0_addr(ram_w32_l1024_id2_0_addr),
    .ram_w32_l1024_id2_0_rdata(ram_w32_l1024_id2_0_rdata),
    .ram_w32_l1024_id2_0_wdata(ram_w32_l1024_id2_0_wdata),
    .ram_w32_l1024_id2_0_wenable(ram_w32_l1024_id2_0_wenable),
    .ram_w32_l1024_id2_0_enable(ram_w32_l1024_id2_0_enable),
    .ram_w32_l1024_id2_1_addr(ram_w32_l1024_id2_1_addr),
    .ram_w32_l1024_id2_1_rdata(ram_w32_l1024_id2_1_rdata),
    .ram_w32_l1024_id2_1_wdata(ram_w32_l1024_id2_1_wdata),
    .ram_w32_l1024_id2_1_wenable(ram_w32_l1024_id2_1_wenable),
    .ram_w32_l1024_id2_1_enable(ram_w32_l1024_id2_1_enable)
  );

  wire [10-1:0] ram_w32_l1024_id3_0_addr;
  wire [32-1:0] ram_w32_l1024_id3_0_rdata;
  wire [32-1:0] ram_w32_l1024_id3_0_wdata;
  wire ram_w32_l1024_id3_0_wenable;
  wire ram_w32_l1024_id3_0_enable;
  wire [10-1:0] ram_w32_l1024_id3_1_addr;
  wire [32-1:0] ram_w32_l1024_id3_1_rdata;
  wire [32-1:0] ram_w32_l1024_id3_1_wdata;
  wire ram_w32_l1024_id3_1_wenable;
  wire ram_w32_l1024_id3_1_enable;
  assign ram_w32_l1024_id3_0_wdata = 'hx;
  assign ram_w32_l1024_id3_0_wenable = 0;

  ram_w32_l1024_id3
  inst_ram_w32_l1024_id3
  (
    .CLK(CLK),
    .ram_w32_l1024_id3_0_addr(ram_w32_l1024_id3_0_addr),
    .ram_w32_l1024_id3_0_rdata(ram_w32_l1024_id3_0_rdata),
    .ram_w32_l1024_id3_0_wdata(ram_w32_l1024_id3_0_wdata),
    .ram_w32_l1024_id3_0_wenable(ram_w32_l1024_id3_0_wenable),
    .ram_w32_l1024_id3_0_enable(ram_w32_l1024_id3_0_enable),
    .ram_w32_l1024_id3_1_addr(ram_w32_l1024_id3_1_addr),
    .ram_w32_l1024_id3_1_rdata(ram_w32_l1024_id3_1_rdata),
    .ram_w32_l1024_id3_1_wdata(ram_w32_l1024_id3_1_wdata),
    .ram_w32_l1024_id3_1_wenable(ram_w32_l1024_id3_1_wenable),
    .ram_w32_l1024_id3_1_enable(ram_w32_l1024_id3_1_enable)
  );

  wire [10-1:0] ram_w32_l1024_id4_0_addr;
  wire [32-1:0] ram_w32_l1024_id4_0_rdata;
  wire [32-1:0] ram_w32_l1024_id4_0_wdata;
  wire ram_w32_l1024_id4_0_wenable;
  wire ram_w32_l1024_id4_0_enable;
  wire [10-1:0] ram_w32_l1024_id4_1_addr;
  wire [32-1:0] ram_w32_l1024_id4_1_rdata;
  wire [32-1:0] ram_w32_l1024_id4_1_wdata;
  wire ram_w32_l1024_id4_1_wenable;
  wire ram_w32_l1024_id4_1_enable;
  assign ram_w32_l1024_id4_0_wdata = 'hx;
  assign ram_w32_l1024_id4_0_wenable = 0;

  ram_w32_l1024_id4
  inst_ram_w32_l1024_id4
  (
    .CLK(CLK),
    .ram_w32_l1024_id4_0_addr(ram_w32_l1024_id4_0_addr),
    .ram_w32_l1024_id4_0_rdata(ram_w32_l1024_id4_0_rdata),
    .ram_w32_l1024_id4_0_wdata(ram_w32_l1024_id4_0_wdata),
    .ram_w32_l1024_id4_0_wenable(ram_w32_l1024_id4_0_wenable),
    .ram_w32_l1024_id4_0_enable(ram_w32_l1024_id4_0_enable),
    .ram_w32_l1024_id4_1_addr(ram_w32_l1024_id4_1_addr),
    .ram_w32_l1024_id4_1_rdata(ram_w32_l1024_id4_1_rdata),
    .ram_w32_l1024_id4_1_wdata(ram_w32_l1024_id4_1_wdata),
    .ram_w32_l1024_id4_1_wenable(ram_w32_l1024_id4_1_wenable),
    .ram_w32_l1024_id4_1_enable(ram_w32_l1024_id4_1_enable)
  );

  wire [10-1:0] ram_w32_l1024_id5_0_addr;
  wire [32-1:0] ram_w32_l1024_id5_0_rdata;
  wire [32-1:0] ram_w32_l1024_id5_0_wdata;
  wire ram_w32_l1024_id5_0_wenable;
  wire ram_w32_l1024_id5_0_enable;
  wire [10-1:0] ram_w32_l1024_id5_1_addr;
  wire [32-1:0] ram_w32_l1024_id5_1_rdata;
  wire [32-1:0] ram_w32_l1024_id5_1_wdata;
  wire ram_w32_l1024_id5_1_wenable;
  wire ram_w32_l1024_id5_1_enable;
  assign ram_w32_l1024_id5_0_wdata = 'hx;
  assign ram_w32_l1024_id5_0_wenable = 0;

  ram_w32_l1024_id5
  inst_ram_w32_l1024_id5
  (
    .CLK(CLK),
    .ram_w32_l1024_id5_0_addr(ram_w32_l1024_id5_0_addr),
    .ram_w32_l1024_id5_0_rdata(ram_w32_l1024_id5_0_rdata),
    .ram_w32_l1024_id5_0_wdata(ram_w32_l1024_id5_0_wdata),
    .ram_w32_l1024_id5_0_wenable(ram_w32_l1024_id5_0_wenable),
    .ram_w32_l1024_id5_0_enable(ram_w32_l1024_id5_0_enable),
    .ram_w32_l1024_id5_1_addr(ram_w32_l1024_id5_1_addr),
    .ram_w32_l1024_id5_1_rdata(ram_w32_l1024_id5_1_rdata),
    .ram_w32_l1024_id5_1_wdata(ram_w32_l1024_id5_1_wdata),
    .ram_w32_l1024_id5_1_wenable(ram_w32_l1024_id5_1_wenable),
    .ram_w32_l1024_id5_1_enable(ram_w32_l1024_id5_1_enable)
  );

  wire [10-1:0] ram_w32_l1024_id6_0_addr;
  wire [32-1:0] ram_w32_l1024_id6_0_rdata;
  wire [32-1:0] ram_w32_l1024_id6_0_wdata;
  wire ram_w32_l1024_id6_0_wenable;
  wire ram_w32_l1024_id6_0_enable;
  wire [10-1:0] ram_w32_l1024_id6_1_addr;
  wire [32-1:0] ram_w32_l1024_id6_1_rdata;
  wire [32-1:0] ram_w32_l1024_id6_1_wdata;
  wire ram_w32_l1024_id6_1_wenable;
  wire ram_w32_l1024_id6_1_enable;
  assign ram_w32_l1024_id6_0_wdata = 'hx;
  assign ram_w32_l1024_id6_0_wenable = 0;

  ram_w32_l1024_id6
  inst_ram_w32_l1024_id6
  (
    .CLK(CLK),
    .ram_w32_l1024_id6_0_addr(ram_w32_l1024_id6_0_addr),
    .ram_w32_l1024_id6_0_rdata(ram_w32_l1024_id6_0_rdata),
    .ram_w32_l1024_id6_0_wdata(ram_w32_l1024_id6_0_wdata),
    .ram_w32_l1024_id6_0_wenable(ram_w32_l1024_id6_0_wenable),
    .ram_w32_l1024_id6_0_enable(ram_w32_l1024_id6_0_enable),
    .ram_w32_l1024_id6_1_addr(ram_w32_l1024_id6_1_addr),
    .ram_w32_l1024_id6_1_rdata(ram_w32_l1024_id6_1_rdata),
    .ram_w32_l1024_id6_1_wdata(ram_w32_l1024_id6_1_wdata),
    .ram_w32_l1024_id6_1_wenable(ram_w32_l1024_id6_1_wenable),
    .ram_w32_l1024_id6_1_enable(ram_w32_l1024_id6_1_enable)
  );

  wire [10-1:0] ram_w32_l1024_id7_0_addr;
  wire [32-1:0] ram_w32_l1024_id7_0_rdata;
  wire [32-1:0] ram_w32_l1024_id7_0_wdata;
  wire ram_w32_l1024_id7_0_wenable;
  wire ram_w32_l1024_id7_0_enable;
  wire [10-1:0] ram_w32_l1024_id7_1_addr;
  wire [32-1:0] ram_w32_l1024_id7_1_rdata;
  wire [32-1:0] ram_w32_l1024_id7_1_wdata;
  wire ram_w32_l1024_id7_1_wenable;
  wire ram_w32_l1024_id7_1_enable;
  assign ram_w32_l1024_id7_0_wdata = 'hx;
  assign ram_w32_l1024_id7_0_wenable = 0;

  ram_w32_l1024_id7
  inst_ram_w32_l1024_id7
  (
    .CLK(CLK),
    .ram_w32_l1024_id7_0_addr(ram_w32_l1024_id7_0_addr),
    .ram_w32_l1024_id7_0_rdata(ram_w32_l1024_id7_0_rdata),
    .ram_w32_l1024_id7_0_wdata(ram_w32_l1024_id7_0_wdata),
    .ram_w32_l1024_id7_0_wenable(ram_w32_l1024_id7_0_wenable),
    .ram_w32_l1024_id7_0_enable(ram_w32_l1024_id7_0_enable),
    .ram_w32_l1024_id7_1_addr(ram_w32_l1024_id7_1_addr),
    .ram_w32_l1024_id7_1_rdata(ram_w32_l1024_id7_1_rdata),
    .ram_w32_l1024_id7_1_wdata(ram_w32_l1024_id7_1_wdata),
    .ram_w32_l1024_id7_1_wenable(ram_w32_l1024_id7_1_wenable),
    .ram_w32_l1024_id7_1_enable(ram_w32_l1024_id7_1_enable)
  );

  wire [10-1:0] ram_w32_l1024_id8_0_addr;
  wire [32-1:0] ram_w32_l1024_id8_0_rdata;
  wire [32-1:0] ram_w32_l1024_id8_0_wdata;
  wire ram_w32_l1024_id8_0_wenable;
  wire ram_w32_l1024_id8_0_enable;
  wire [10-1:0] ram_w32_l1024_id8_1_addr;
  wire [32-1:0] ram_w32_l1024_id8_1_rdata;
  wire [32-1:0] ram_w32_l1024_id8_1_wdata;
  wire ram_w32_l1024_id8_1_wenable;
  wire ram_w32_l1024_id8_1_enable;
  assign ram_w32_l1024_id8_0_wdata = 'hx;
  assign ram_w32_l1024_id8_0_wenable = 0;

  ram_w32_l1024_id8
  inst_ram_w32_l1024_id8
  (
    .CLK(CLK),
    .ram_w32_l1024_id8_0_addr(ram_w32_l1024_id8_0_addr),
    .ram_w32_l1024_id8_0_rdata(ram_w32_l1024_id8_0_rdata),
    .ram_w32_l1024_id8_0_wdata(ram_w32_l1024_id8_0_wdata),
    .ram_w32_l1024_id8_0_wenable(ram_w32_l1024_id8_0_wenable),
    .ram_w32_l1024_id8_0_enable(ram_w32_l1024_id8_0_enable),
    .ram_w32_l1024_id8_1_addr(ram_w32_l1024_id8_1_addr),
    .ram_w32_l1024_id8_1_rdata(ram_w32_l1024_id8_1_rdata),
    .ram_w32_l1024_id8_1_wdata(ram_w32_l1024_id8_1_wdata),
    .ram_w32_l1024_id8_1_wenable(ram_w32_l1024_id8_1_wenable),
    .ram_w32_l1024_id8_1_enable(ram_w32_l1024_id8_1_enable)
  );

  wire [10-1:0] ram_w32_l1024_id9_0_addr;
  wire [32-1:0] ram_w32_l1024_id9_0_rdata;
  wire [32-1:0] ram_w32_l1024_id9_0_wdata;
  wire ram_w32_l1024_id9_0_wenable;
  wire ram_w32_l1024_id9_0_enable;
  wire [10-1:0] ram_w32_l1024_id9_1_addr;
  wire [32-1:0] ram_w32_l1024_id9_1_rdata;
  wire [32-1:0] ram_w32_l1024_id9_1_wdata;
  wire ram_w32_l1024_id9_1_wenable;
  wire ram_w32_l1024_id9_1_enable;
  assign ram_w32_l1024_id9_0_wdata = 'hx;
  assign ram_w32_l1024_id9_0_wenable = 0;

  ram_w32_l1024_id9
  inst_ram_w32_l1024_id9
  (
    .CLK(CLK),
    .ram_w32_l1024_id9_0_addr(ram_w32_l1024_id9_0_addr),
    .ram_w32_l1024_id9_0_rdata(ram_w32_l1024_id9_0_rdata),
    .ram_w32_l1024_id9_0_wdata(ram_w32_l1024_id9_0_wdata),
    .ram_w32_l1024_id9_0_wenable(ram_w32_l1024_id9_0_wenable),
    .ram_w32_l1024_id9_0_enable(ram_w32_l1024_id9_0_enable),
    .ram_w32_l1024_id9_1_addr(ram_w32_l1024_id9_1_addr),
    .ram_w32_l1024_id9_1_rdata(ram_w32_l1024_id9_1_rdata),
    .ram_w32_l1024_id9_1_wdata(ram_w32_l1024_id9_1_wdata),
    .ram_w32_l1024_id9_1_wenable(ram_w32_l1024_id9_1_wenable),
    .ram_w32_l1024_id9_1_enable(ram_w32_l1024_id9_1_enable)
  );

  wire [10-1:0] ram_w32_l1024_id10_0_addr;
  wire [32-1:0] ram_w32_l1024_id10_0_rdata;
  wire [32-1:0] ram_w32_l1024_id10_0_wdata;
  wire ram_w32_l1024_id10_0_wenable;
  wire ram_w32_l1024_id10_0_enable;
  wire [10-1:0] ram_w32_l1024_id10_1_addr;
  wire [32-1:0] ram_w32_l1024_id10_1_rdata;
  wire [32-1:0] ram_w32_l1024_id10_1_wdata;
  wire ram_w32_l1024_id10_1_wenable;
  wire ram_w32_l1024_id10_1_enable;
  assign ram_w32_l1024_id10_0_wdata = 'hx;
  assign ram_w32_l1024_id10_0_wenable = 0;

  ram_w32_l1024_id10
  inst_ram_w32_l1024_id10
  (
    .CLK(CLK),
    .ram_w32_l1024_id10_0_addr(ram_w32_l1024_id10_0_addr),
    .ram_w32_l1024_id10_0_rdata(ram_w32_l1024_id10_0_rdata),
    .ram_w32_l1024_id10_0_wdata(ram_w32_l1024_id10_0_wdata),
    .ram_w32_l1024_id10_0_wenable(ram_w32_l1024_id10_0_wenable),
    .ram_w32_l1024_id10_0_enable(ram_w32_l1024_id10_0_enable),
    .ram_w32_l1024_id10_1_addr(ram_w32_l1024_id10_1_addr),
    .ram_w32_l1024_id10_1_rdata(ram_w32_l1024_id10_1_rdata),
    .ram_w32_l1024_id10_1_wdata(ram_w32_l1024_id10_1_wdata),
    .ram_w32_l1024_id10_1_wenable(ram_w32_l1024_id10_1_wenable),
    .ram_w32_l1024_id10_1_enable(ram_w32_l1024_id10_1_enable)
  );

  wire [9-1:0] cparam_conv2d_25_act_num_col;
  wire [9-1:0] cparam_conv2d_25_act_num_row;
  wire [11-1:0] cparam_conv2d_25_filter_num_och;
  wire [1-1:0] cparam_conv2d_25_bias_scala;
  wire [11-1:0] cparam_conv2d_25_bias_num;
  wire [1-1:0] cparam_conv2d_25_scale_scala;
  wire [1-1:0] cparam_conv2d_25_scale_num;
  wire [1-1:0] cparam_conv2d_25_vshamt_mul_scala;
  wire [1-1:0] cparam_conv2d_25_vshamt_mul_num;
  wire [1-1:0] cparam_conv2d_25_vshamt_sum_scala;
  wire [1-1:0] cparam_conv2d_25_vshamt_sum_num;
  wire [1-1:0] cparam_conv2d_25_vshamt_out_scala;
  wire [1-1:0] cparam_conv2d_25_vshamt_out_num;
  wire [1-1:0] cparam_conv2d_25_cshamt_mul_value;
  wire [1-1:0] cparam_conv2d_25_cshamt_sum_value;
  wire [5-1:0] cparam_conv2d_25_cshamt_out_value;
  wire [1-1:0] cparam_conv2d_25_act_func_index;
  wire [9-1:0] cparam_conv2d_25_out_num_col;
  wire [9-1:0] cparam_conv2d_25_out_num_row;
  wire [1-1:0] cparam_conv2d_25_pad_col_left;
  wire [1-1:0] cparam_conv2d_25_pad_row_top;
  wire [9-1:0] cparam_conv2d_25_max_col_count;
  wire [9-1:0] cparam_conv2d_25_max_row_count;
  wire [1-1:0] cparam_conv2d_25_max_bat_count;
  wire [10-1:0] cparam_conv2d_25_max_och_count;
  wire [4-1:0] cparam_conv2d_25_och_count_step;
  wire [1-1:0] cparam_conv2d_25_dma_flag_conds_0;
  wire [1-1:0] cparam_conv2d_25_dma_flag_conds_1;
  wire [1-1:0] cparam_conv2d_25_dma_flag_conds_2;
  wire signed [32-1:0] cparam_conv2d_25_act_offset_values_0;
  wire signed [32-1:0] cparam_conv2d_25_act_offset_values_1;
  wire signed [32-1:0] cparam_conv2d_25_act_offset_values_2;
  wire [15-1:0] cparam_conv2d_25_act_row_step;
  wire [22-1:0] cparam_conv2d_25_act_bat_step;
  wire [13-1:0] cparam_conv2d_25_act_read_size;
  wire [10-1:0] cparam_conv2d_25_act_read_block;
  wire [12-1:0] cparam_conv2d_25_act_read_step;
  wire [15-1:0] cparam_conv2d_25_filter_base_step;
  wire [13-1:0] cparam_conv2d_25_filter_read_size;
  wire [10-1:0] cparam_conv2d_25_filter_read_block;
  wire [10-1:0] cparam_conv2d_25_filter_read_step;
  wire [1-1:0] cparam_conv2d_25_out_offset_values_0;
  wire [13-1:0] cparam_conv2d_25_out_col_step;
  wire [16-1:0] cparam_conv2d_25_out_row_step;
  wire [24-1:0] cparam_conv2d_25_out_bat_step;
  wire [6-1:0] cparam_conv2d_25_out_och_step;
  wire [4-1:0] cparam_conv2d_25_out_write_size;
  wire [4-1:0] cparam_conv2d_25_out_write_size_res;
  wire [1-1:0] cparam_conv2d_25_out_write_block;
  wire [1-1:0] cparam_conv2d_25_keep_filter;
  wire [1-1:0] cparam_conv2d_25_keep_input;
  wire [1-1:0] cparam_conv2d_25_data_stationary;
  wire [4-1:0] cparam_conv2d_25_stream_num_ops;
  wire [4-1:0] cparam_conv2d_25_stream_num_ops_res;
  wire [4-1:0] cparam_conv2d_25_stream_num_ops_par;
  wire [4-1:0] cparam_conv2d_25_stream_num_ops_res_par;
  wire [10-1:0] cparam_conv2d_25_stream_reduce_size;
  wire [10-1:0] cparam_conv2d_25_stream_aligned_reduce_size;
  wire [1-1:0] cparam_conv2d_25_stream_omit_mask;
  wire [2-1:0] cparam_conv2d_25_col_select_initval;
  wire [1-1:0] cparam_conv2d_25_stride_col_par_col;
  wire [1-1:0] cparam_conv2d_25_stride_row_par_row;
  wire [1-1:0] cparam_conv2d_25_stride_col_mod_filter_num;
  wire [2-1:0] cparam_conv2d_25_filter_num_col_minus_stride_col_mod;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_0;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_1;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_2;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_3;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_4;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_5;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_6;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_7;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_8;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_9;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_10;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_11;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_12;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_13;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_14;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_15;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_16;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_17;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_18;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_19;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_20;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_21;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_22;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_23;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_24;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_25;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_conds_26;
  wire [1-1:0] cparam_conv2d_25_inc_act_laddr_small;
  wire [10-1:0] cparam_conv2d_25_inc_act_laddr_large;
  wire [11-1:0] cparam_conv2d_25_inc_out_laddr_col;
  wire [1-1:0] cparam_conv2d_25_stream_act_local_small_offset;
  wire signed [11-1:0] cparam_conv2d_25_stream_act_local_large_offset;
  wire [1-1:0] cparam_conv2d_25_stream_act_local_small_flags_0;
  wire [1-1:0] cparam_conv2d_25_stream_act_local_small_flags_1;
  wire [1-1:0] cparam_conv2d_25_stream_act_local_small_flags_2;
  wire [1-1:0] cparam_conv2d_25_stream_act_local_large_flags_0;
  wire [1-1:0] cparam_conv2d_25_stream_act_local_large_flags_1;
  wire [1-1:0] cparam_conv2d_25_stream_act_local_large_flags_2;
  wire [1-1:0] cparam_conv2d_25_inc_sync_out;
  wire [1-1:0] cparam_conv2d_25_inc_sync_out_res;
  reg [3-1:0] conv2d_25_control_param_index;
  assign cparam_conv2d_25_act_num_col = (conv2d_25_control_param_index == 0)? 32'h1a0 : 
                                        (conv2d_25_control_param_index == 1)? 32'hd0 : 
                                        (conv2d_25_control_param_index == 2)? 32'h68 : 
                                        (conv2d_25_control_param_index == 3)? 32'h34 : 
                                        (conv2d_25_control_param_index == 4)? 32'h1a : 
                                        (conv2d_25_control_param_index == 5)? 32'hd : 32'hc;
  assign cparam_conv2d_25_act_num_row = (conv2d_25_control_param_index == 0)? 32'h1a0 : 
                                        (conv2d_25_control_param_index == 1)? 32'hd0 : 
                                        (conv2d_25_control_param_index == 2)? 32'h68 : 
                                        (conv2d_25_control_param_index == 3)? 32'h34 : 
                                        (conv2d_25_control_param_index == 4)? 32'h1a : 
                                        (conv2d_25_control_param_index == 5)? 32'hd : 32'hc;
  assign cparam_conv2d_25_filter_num_och = (conv2d_25_control_param_index == 0)? 32'h10 : 
                                           (conv2d_25_control_param_index == 1)? 32'h20 : 
                                           (conv2d_25_control_param_index == 2)? 32'h40 : 
                                           (conv2d_25_control_param_index == 3)? 32'h80 : 
                                           (conv2d_25_control_param_index == 4)? 32'h100 : 
                                           (conv2d_25_control_param_index == 5)? 32'h200 : 32'h400;
  assign cparam_conv2d_25_bias_scala = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                       (conv2d_25_control_param_index == 1)? 32'h0 : 
                                       (conv2d_25_control_param_index == 2)? 32'h0 : 
                                       (conv2d_25_control_param_index == 3)? 32'h0 : 
                                       (conv2d_25_control_param_index == 4)? 32'h0 : 
                                       (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_bias_num = (conv2d_25_control_param_index == 0)? 32'h10 : 
                                     (conv2d_25_control_param_index == 1)? 32'h20 : 
                                     (conv2d_25_control_param_index == 2)? 32'h40 : 
                                     (conv2d_25_control_param_index == 3)? 32'h80 : 
                                     (conv2d_25_control_param_index == 4)? 32'h100 : 
                                     (conv2d_25_control_param_index == 5)? 32'h200 : 32'h400;
  assign cparam_conv2d_25_scale_scala = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                        (conv2d_25_control_param_index == 1)? 32'h1 : 
                                        (conv2d_25_control_param_index == 2)? 32'h1 : 
                                        (conv2d_25_control_param_index == 3)? 32'h1 : 
                                        (conv2d_25_control_param_index == 4)? 32'h1 : 
                                        (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_scale_num = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                      (conv2d_25_control_param_index == 1)? 32'h1 : 
                                      (conv2d_25_control_param_index == 2)? 32'h1 : 
                                      (conv2d_25_control_param_index == 3)? 32'h1 : 
                                      (conv2d_25_control_param_index == 4)? 32'h1 : 
                                      (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_vshamt_mul_scala = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                             (conv2d_25_control_param_index == 1)? 32'h0 : 
                                             (conv2d_25_control_param_index == 2)? 32'h0 : 
                                             (conv2d_25_control_param_index == 3)? 32'h0 : 
                                             (conv2d_25_control_param_index == 4)? 32'h0 : 
                                             (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_vshamt_mul_num = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                           (conv2d_25_control_param_index == 1)? 32'h0 : 
                                           (conv2d_25_control_param_index == 2)? 32'h0 : 
                                           (conv2d_25_control_param_index == 3)? 32'h0 : 
                                           (conv2d_25_control_param_index == 4)? 32'h0 : 
                                           (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_vshamt_sum_scala = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                             (conv2d_25_control_param_index == 1)? 32'h0 : 
                                             (conv2d_25_control_param_index == 2)? 32'h0 : 
                                             (conv2d_25_control_param_index == 3)? 32'h0 : 
                                             (conv2d_25_control_param_index == 4)? 32'h0 : 
                                             (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_vshamt_sum_num = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                           (conv2d_25_control_param_index == 1)? 32'h0 : 
                                           (conv2d_25_control_param_index == 2)? 32'h0 : 
                                           (conv2d_25_control_param_index == 3)? 32'h0 : 
                                           (conv2d_25_control_param_index == 4)? 32'h0 : 
                                           (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_vshamt_out_scala = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                             (conv2d_25_control_param_index == 1)? 32'h0 : 
                                             (conv2d_25_control_param_index == 2)? 32'h0 : 
                                             (conv2d_25_control_param_index == 3)? 32'h0 : 
                                             (conv2d_25_control_param_index == 4)? 32'h0 : 
                                             (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_vshamt_out_num = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                           (conv2d_25_control_param_index == 1)? 32'h0 : 
                                           (conv2d_25_control_param_index == 2)? 32'h0 : 
                                           (conv2d_25_control_param_index == 3)? 32'h0 : 
                                           (conv2d_25_control_param_index == 4)? 32'h0 : 
                                           (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_cshamt_mul_value = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                             (conv2d_25_control_param_index == 1)? 32'h0 : 
                                             (conv2d_25_control_param_index == 2)? 32'h0 : 
                                             (conv2d_25_control_param_index == 3)? 32'h0 : 
                                             (conv2d_25_control_param_index == 4)? 32'h0 : 
                                             (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_cshamt_sum_value = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                             (conv2d_25_control_param_index == 1)? 32'h0 : 
                                             (conv2d_25_control_param_index == 2)? 32'h0 : 
                                             (conv2d_25_control_param_index == 3)? 32'h0 : 
                                             (conv2d_25_control_param_index == 4)? 32'h0 : 
                                             (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_cshamt_out_value = (conv2d_25_control_param_index == 0)? 32'h1e : 
                                             (conv2d_25_control_param_index == 1)? 32'h1d : 
                                             (conv2d_25_control_param_index == 2)? 32'h1c : 
                                             (conv2d_25_control_param_index == 3)? 32'h1c : 
                                             (conv2d_25_control_param_index == 4)? 32'h1b : 
                                             (conv2d_25_control_param_index == 5)? 32'h1b : 32'h1b;
  assign cparam_conv2d_25_act_func_index = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                           (conv2d_25_control_param_index == 1)? 32'h0 : 
                                           (conv2d_25_control_param_index == 2)? 32'h0 : 
                                           (conv2d_25_control_param_index == 3)? 32'h0 : 
                                           (conv2d_25_control_param_index == 4)? 32'h0 : 
                                           (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_out_num_col = (conv2d_25_control_param_index == 0)? 32'h1a0 : 
                                        (conv2d_25_control_param_index == 1)? 32'hd0 : 
                                        (conv2d_25_control_param_index == 2)? 32'h68 : 
                                        (conv2d_25_control_param_index == 3)? 32'h34 : 
                                        (conv2d_25_control_param_index == 4)? 32'h1a : 
                                        (conv2d_25_control_param_index == 5)? 32'hd : 32'hc;
  assign cparam_conv2d_25_out_num_row = (conv2d_25_control_param_index == 0)? 32'h1a0 : 
                                        (conv2d_25_control_param_index == 1)? 32'hd0 : 
                                        (conv2d_25_control_param_index == 2)? 32'h68 : 
                                        (conv2d_25_control_param_index == 3)? 32'h34 : 
                                        (conv2d_25_control_param_index == 4)? 32'h1a : 
                                        (conv2d_25_control_param_index == 5)? 32'hd : 32'hc;
  assign cparam_conv2d_25_pad_col_left = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                         (conv2d_25_control_param_index == 1)? 32'h1 : 
                                         (conv2d_25_control_param_index == 2)? 32'h1 : 
                                         (conv2d_25_control_param_index == 3)? 32'h1 : 
                                         (conv2d_25_control_param_index == 4)? 32'h1 : 
                                         (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_pad_row_top = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                        (conv2d_25_control_param_index == 1)? 32'h1 : 
                                        (conv2d_25_control_param_index == 2)? 32'h1 : 
                                        (conv2d_25_control_param_index == 3)? 32'h1 : 
                                        (conv2d_25_control_param_index == 4)? 32'h1 : 
                                        (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_max_col_count = (conv2d_25_control_param_index == 0)? 32'h19f : 
                                          (conv2d_25_control_param_index == 1)? 32'hcf : 
                                          (conv2d_25_control_param_index == 2)? 32'h67 : 
                                          (conv2d_25_control_param_index == 3)? 32'h33 : 
                                          (conv2d_25_control_param_index == 4)? 32'h19 : 
                                          (conv2d_25_control_param_index == 5)? 32'hc : 32'hb;
  assign cparam_conv2d_25_max_row_count = (conv2d_25_control_param_index == 0)? 32'h19f : 
                                          (conv2d_25_control_param_index == 1)? 32'hcf : 
                                          (conv2d_25_control_param_index == 2)? 32'h67 : 
                                          (conv2d_25_control_param_index == 3)? 32'h33 : 
                                          (conv2d_25_control_param_index == 4)? 32'h19 : 
                                          (conv2d_25_control_param_index == 5)? 32'hc : 32'hb;
  assign cparam_conv2d_25_max_bat_count = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                          (conv2d_25_control_param_index == 1)? 32'h0 : 
                                          (conv2d_25_control_param_index == 2)? 32'h0 : 
                                          (conv2d_25_control_param_index == 3)? 32'h0 : 
                                          (conv2d_25_control_param_index == 4)? 32'h0 : 
                                          (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_max_och_count = (conv2d_25_control_param_index == 0)? 32'hf : 
                                          (conv2d_25_control_param_index == 1)? 32'h1e : 
                                          (conv2d_25_control_param_index == 2)? 32'h3c : 
                                          (conv2d_25_control_param_index == 3)? 32'h78 : 
                                          (conv2d_25_control_param_index == 4)? 32'hfc : 
                                          (conv2d_25_control_param_index == 5)? 32'h1fe : 32'h3ff;
  assign cparam_conv2d_25_och_count_step = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                           (conv2d_25_control_param_index == 1)? 32'h2 : 
                                           (conv2d_25_control_param_index == 2)? 32'h4 : 
                                           (conv2d_25_control_param_index == 3)? 32'h8 : 
                                           (conv2d_25_control_param_index == 4)? 32'h4 : 
                                           (conv2d_25_control_param_index == 5)? 32'h2 : 32'h1;
  assign cparam_conv2d_25_dma_flag_conds_0 = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                             (conv2d_25_control_param_index == 1)? 32'h1 : 
                                             (conv2d_25_control_param_index == 2)? 32'h1 : 
                                             (conv2d_25_control_param_index == 3)? 32'h1 : 
                                             (conv2d_25_control_param_index == 4)? 32'h1 : 
                                             (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_dma_flag_conds_1 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                             (conv2d_25_control_param_index == 1)? 32'h0 : 
                                             (conv2d_25_control_param_index == 2)? 32'h0 : 
                                             (conv2d_25_control_param_index == 3)? 32'h0 : 
                                             (conv2d_25_control_param_index == 4)? 32'h0 : 
                                             (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_dma_flag_conds_2 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                             (conv2d_25_control_param_index == 1)? 32'h0 : 
                                             (conv2d_25_control_param_index == 2)? 32'h0 : 
                                             (conv2d_25_control_param_index == 3)? 32'h0 : 
                                             (conv2d_25_control_param_index == 4)? 32'h0 : 
                                             (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_act_offset_values_0 = (conv2d_25_control_param_index == 0)? -32'sh1380 : 
                                                (conv2d_25_control_param_index == 1)? -32'sh3400 : 
                                                (conv2d_25_control_param_index == 2)? -32'sh3400 : 
                                                (conv2d_25_control_param_index == 3)? -32'sh3400 : 
                                                (conv2d_25_control_param_index == 4)? -32'sh3400 : 
                                                (conv2d_25_control_param_index == 5)? -32'sh3400 : -32'sh6000;
  assign cparam_conv2d_25_act_offset_values_1 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_act_offset_values_2 = (conv2d_25_control_param_index == 0)? 32'h1380 : 
                                                (conv2d_25_control_param_index == 1)? 32'h3400 : 
                                                (conv2d_25_control_param_index == 2)? 32'h3400 : 
                                                (conv2d_25_control_param_index == 3)? 32'h3400 : 
                                                (conv2d_25_control_param_index == 4)? 32'h3400 : 
                                                (conv2d_25_control_param_index == 5)? 32'h3400 : 32'h6000;
  assign cparam_conv2d_25_act_row_step = (conv2d_25_control_param_index == 0)? 32'h1380 : 
                                         (conv2d_25_control_param_index == 1)? 32'h3400 : 
                                         (conv2d_25_control_param_index == 2)? 32'h3400 : 
                                         (conv2d_25_control_param_index == 3)? 32'h3400 : 
                                         (conv2d_25_control_param_index == 4)? 32'h3400 : 
                                         (conv2d_25_control_param_index == 5)? 32'h3400 : 32'h6000;
  assign cparam_conv2d_25_act_bat_step = (conv2d_25_control_param_index == 0)? 32'h1fb000 : 
                                         (conv2d_25_control_param_index == 1)? 32'h2a4000 : 
                                         (conv2d_25_control_param_index == 2)? 32'h152000 : 
                                         (conv2d_25_control_param_index == 3)? 32'ha9000 : 
                                         (conv2d_25_control_param_index == 4)? 32'h54800 : 
                                         (conv2d_25_control_param_index == 5)? 32'h2a400 : 32'h48000;
  assign cparam_conv2d_25_act_read_size = (conv2d_25_control_param_index == 0)? 32'h4e0 : 
                                          (conv2d_25_control_param_index == 1)? 32'hd00 : 
                                          (conv2d_25_control_param_index == 2)? 32'hd00 : 
                                          (conv2d_25_control_param_index == 3)? 32'hd00 : 
                                          (conv2d_25_control_param_index == 4)? 32'hd00 : 
                                          (conv2d_25_control_param_index == 5)? 32'hd00 : 32'h1800;
  assign cparam_conv2d_25_act_read_block = (conv2d_25_control_param_index == 0)? 32'h3 : 
                                           (conv2d_25_control_param_index == 1)? 32'h10 : 
                                           (conv2d_25_control_param_index == 2)? 32'h20 : 
                                           (conv2d_25_control_param_index == 3)? 32'h40 : 
                                           (conv2d_25_control_param_index == 4)? 32'h80 : 
                                           (conv2d_25_control_param_index == 5)? 32'h100 : 32'h200;
  assign cparam_conv2d_25_act_read_step = (conv2d_25_control_param_index == 0)? 32'h1a1 : 
                                          (conv2d_25_control_param_index == 1)? 32'h460 : 
                                          (conv2d_25_control_param_index == 2)? 32'h460 : 
                                          (conv2d_25_control_param_index == 3)? 32'h480 : 
                                          (conv2d_25_control_param_index == 4)? 32'h480 : 
                                          (conv2d_25_control_param_index == 5)? 32'h500 : 32'h800;
  assign cparam_conv2d_25_filter_base_step = (conv2d_25_control_param_index == 0)? 32'h6c : 
                                             (conv2d_25_control_param_index == 1)? 32'h480 : 
                                             (conv2d_25_control_param_index == 2)? 32'h1200 : 
                                             (conv2d_25_control_param_index == 3)? 32'h4800 : 
                                             (conv2d_25_control_param_index == 4)? 32'h4800 : 
                                             (conv2d_25_control_param_index == 5)? 32'h4800 : 32'h4800;
  assign cparam_conv2d_25_filter_read_size = (conv2d_25_control_param_index == 0)? 32'h1b : 
                                             (conv2d_25_control_param_index == 1)? 32'h120 : 
                                             (conv2d_25_control_param_index == 2)? 32'h480 : 
                                             (conv2d_25_control_param_index == 3)? 32'h1200 : 
                                             (conv2d_25_control_param_index == 4)? 32'h1200 : 
                                             (conv2d_25_control_param_index == 5)? 32'h1200 : 32'h1200;
  assign cparam_conv2d_25_filter_read_block = (conv2d_25_control_param_index == 0)? 32'h3 : 
                                              (conv2d_25_control_param_index == 1)? 32'h10 : 
                                              (conv2d_25_control_param_index == 2)? 32'h20 : 
                                              (conv2d_25_control_param_index == 3)? 32'h40 : 
                                              (conv2d_25_control_param_index == 4)? 32'h80 : 
                                              (conv2d_25_control_param_index == 5)? 32'h100 : 32'h200;
  assign cparam_conv2d_25_filter_read_step = (conv2d_25_control_param_index == 0)? 32'h3 : 
                                             (conv2d_25_control_param_index == 1)? 32'h20 : 
                                             (conv2d_25_control_param_index == 2)? 32'h80 : 
                                             (conv2d_25_control_param_index == 3)? 32'h200 : 
                                             (conv2d_25_control_param_index == 4)? 32'h200 : 
                                             (conv2d_25_control_param_index == 5)? 32'h200 : 32'h200;
  assign cparam_conv2d_25_out_offset_values_0 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_out_col_step = (conv2d_25_control_param_index == 0)? 32'h40 : 
                                         (conv2d_25_control_param_index == 1)? 32'h80 : 
                                         (conv2d_25_control_param_index == 2)? 32'h100 : 
                                         (conv2d_25_control_param_index == 3)? 32'h200 : 
                                         (conv2d_25_control_param_index == 4)? 32'h400 : 
                                         (conv2d_25_control_param_index == 5)? 32'h800 : 32'h1000;
  assign cparam_conv2d_25_out_row_step = (conv2d_25_control_param_index == 0)? 32'h6800 : 
                                         (conv2d_25_control_param_index == 1)? 32'h6800 : 
                                         (conv2d_25_control_param_index == 2)? 32'h6800 : 
                                         (conv2d_25_control_param_index == 3)? 32'h6800 : 
                                         (conv2d_25_control_param_index == 4)? 32'h6800 : 
                                         (conv2d_25_control_param_index == 5)? 32'h6800 : 32'hc000;
  assign cparam_conv2d_25_out_bat_step = (conv2d_25_control_param_index == 0)? 32'ha90000 : 
                                         (conv2d_25_control_param_index == 1)? 32'h548000 : 
                                         (conv2d_25_control_param_index == 2)? 32'h2a4000 : 
                                         (conv2d_25_control_param_index == 3)? 32'h152000 : 
                                         (conv2d_25_control_param_index == 4)? 32'ha9000 : 
                                         (conv2d_25_control_param_index == 5)? 32'h54800 : 32'h90000;
  assign cparam_conv2d_25_out_och_step = (conv2d_25_control_param_index == 0)? 32'h4 : 
                                         (conv2d_25_control_param_index == 1)? 32'h8 : 
                                         (conv2d_25_control_param_index == 2)? 32'h10 : 
                                         (conv2d_25_control_param_index == 3)? 32'h20 : 
                                         (conv2d_25_control_param_index == 4)? 32'h10 : 
                                         (conv2d_25_control_param_index == 5)? 32'h8 : 32'h4;
  assign cparam_conv2d_25_out_write_size = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                           (conv2d_25_control_param_index == 1)? 32'h2 : 
                                           (conv2d_25_control_param_index == 2)? 32'h4 : 
                                           (conv2d_25_control_param_index == 3)? 32'h8 : 
                                           (conv2d_25_control_param_index == 4)? 32'h4 : 
                                           (conv2d_25_control_param_index == 5)? 32'h2 : 32'h1;
  assign cparam_conv2d_25_out_write_size_res = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                               (conv2d_25_control_param_index == 1)? 32'h2 : 
                                               (conv2d_25_control_param_index == 2)? 32'h4 : 
                                               (conv2d_25_control_param_index == 3)? 32'h8 : 
                                               (conv2d_25_control_param_index == 4)? 32'h4 : 
                                               (conv2d_25_control_param_index == 5)? 32'h2 : 32'h1;
  assign cparam_conv2d_25_out_write_block = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                            (conv2d_25_control_param_index == 1)? 32'h0 : 
                                            (conv2d_25_control_param_index == 2)? 32'h0 : 
                                            (conv2d_25_control_param_index == 3)? 32'h0 : 
                                            (conv2d_25_control_param_index == 4)? 32'h0 : 
                                            (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_keep_filter = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                        (conv2d_25_control_param_index == 1)? 32'h0 : 
                                        (conv2d_25_control_param_index == 2)? 32'h0 : 
                                        (conv2d_25_control_param_index == 3)? 32'h0 : 
                                        (conv2d_25_control_param_index == 4)? 32'h0 : 
                                        (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_keep_input = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                       (conv2d_25_control_param_index == 1)? 32'h0 : 
                                       (conv2d_25_control_param_index == 2)? 32'h0 : 
                                       (conv2d_25_control_param_index == 3)? 32'h0 : 
                                       (conv2d_25_control_param_index == 4)? 32'h0 : 
                                       (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_data_stationary = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                            (conv2d_25_control_param_index == 1)? 32'h0 : 
                                            (conv2d_25_control_param_index == 2)? 32'h0 : 
                                            (conv2d_25_control_param_index == 3)? 32'h0 : 
                                            (conv2d_25_control_param_index == 4)? 32'h0 : 
                                            (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_stream_num_ops = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                           (conv2d_25_control_param_index == 1)? 32'h2 : 
                                           (conv2d_25_control_param_index == 2)? 32'h4 : 
                                           (conv2d_25_control_param_index == 3)? 32'h8 : 
                                           (conv2d_25_control_param_index == 4)? 32'h4 : 
                                           (conv2d_25_control_param_index == 5)? 32'h2 : 32'h1;
  assign cparam_conv2d_25_stream_num_ops_res = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                               (conv2d_25_control_param_index == 1)? 32'h2 : 
                                               (conv2d_25_control_param_index == 2)? 32'h4 : 
                                               (conv2d_25_control_param_index == 3)? 32'h8 : 
                                               (conv2d_25_control_param_index == 4)? 32'h4 : 
                                               (conv2d_25_control_param_index == 5)? 32'h2 : 32'h1;
  assign cparam_conv2d_25_stream_num_ops_par = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                               (conv2d_25_control_param_index == 1)? 32'h2 : 
                                               (conv2d_25_control_param_index == 2)? 32'h4 : 
                                               (conv2d_25_control_param_index == 3)? 32'h8 : 
                                               (conv2d_25_control_param_index == 4)? 32'h4 : 
                                               (conv2d_25_control_param_index == 5)? 32'h2 : 32'h1;
  assign cparam_conv2d_25_stream_num_ops_res_par = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h2 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h4 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h8 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h4 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h2 : 32'h1;
  assign cparam_conv2d_25_stream_reduce_size = (conv2d_25_control_param_index == 0)? 32'h3 : 
                                               (conv2d_25_control_param_index == 1)? 32'h10 : 
                                               (conv2d_25_control_param_index == 2)? 32'h20 : 
                                               (conv2d_25_control_param_index == 3)? 32'h40 : 
                                               (conv2d_25_control_param_index == 4)? 32'h80 : 
                                               (conv2d_25_control_param_index == 5)? 32'h100 : 32'h200;
  assign cparam_conv2d_25_stream_aligned_reduce_size = (conv2d_25_control_param_index == 0)? 32'h3 : 
                                                       (conv2d_25_control_param_index == 1)? 32'h10 : 
                                                       (conv2d_25_control_param_index == 2)? 32'h20 : 
                                                       (conv2d_25_control_param_index == 3)? 32'h40 : 
                                                       (conv2d_25_control_param_index == 4)? 32'h80 : 
                                                       (conv2d_25_control_param_index == 5)? 32'h100 : 32'h200;
  assign cparam_conv2d_25_stream_omit_mask = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                             (conv2d_25_control_param_index == 1)? 32'h0 : 
                                             (conv2d_25_control_param_index == 2)? 32'h0 : 
                                             (conv2d_25_control_param_index == 3)? 32'h0 : 
                                             (conv2d_25_control_param_index == 4)? 32'h0 : 
                                             (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_col_select_initval = (conv2d_25_control_param_index == 0)? 32'h2 : 
                                               (conv2d_25_control_param_index == 1)? 32'h2 : 
                                               (conv2d_25_control_param_index == 2)? 32'h2 : 
                                               (conv2d_25_control_param_index == 3)? 32'h2 : 
                                               (conv2d_25_control_param_index == 4)? 32'h2 : 
                                               (conv2d_25_control_param_index == 5)? 32'h2 : 32'h2;
  assign cparam_conv2d_25_stride_col_par_col = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                               (conv2d_25_control_param_index == 1)? 32'h1 : 
                                               (conv2d_25_control_param_index == 2)? 32'h1 : 
                                               (conv2d_25_control_param_index == 3)? 32'h1 : 
                                               (conv2d_25_control_param_index == 4)? 32'h1 : 
                                               (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_stride_row_par_row = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                               (conv2d_25_control_param_index == 1)? 32'h1 : 
                                               (conv2d_25_control_param_index == 2)? 32'h1 : 
                                               (conv2d_25_control_param_index == 3)? 32'h1 : 
                                               (conv2d_25_control_param_index == 4)? 32'h1 : 
                                               (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_stride_col_mod_filter_num = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                                      (conv2d_25_control_param_index == 1)? 32'h1 : 
                                                      (conv2d_25_control_param_index == 2)? 32'h1 : 
                                                      (conv2d_25_control_param_index == 3)? 32'h1 : 
                                                      (conv2d_25_control_param_index == 4)? 32'h1 : 
                                                      (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_filter_num_col_minus_stride_col_mod = (conv2d_25_control_param_index == 0)? 32'h2 : 
                                                                (conv2d_25_control_param_index == 1)? 32'h2 : 
                                                                (conv2d_25_control_param_index == 2)? 32'h2 : 
                                                                (conv2d_25_control_param_index == 3)? 32'h2 : 
                                                                (conv2d_25_control_param_index == 4)? 32'h2 : 
                                                                (conv2d_25_control_param_index == 5)? 32'h2 : 32'h2;
  assign cparam_conv2d_25_inc_act_laddr_conds_0 = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 1)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 2)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 3)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 4)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_inc_act_laddr_conds_1 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_2 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_3 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_4 = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 1)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 2)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 3)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 4)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_inc_act_laddr_conds_5 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_6 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_7 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                  (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_8 = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 1)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 2)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 3)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 4)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_inc_act_laddr_conds_9 = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 1)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 2)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 3)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 4)? 32'h1 : 
                                                  (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_inc_act_laddr_conds_10 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_11 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_12 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_13 = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_inc_act_laddr_conds_14 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_15 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_16 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_17 = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_inc_act_laddr_conds_18 = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_inc_act_laddr_conds_19 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_20 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_21 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_22 = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_inc_act_laddr_conds_23 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_24 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_25 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_conds_26 = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 1)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 2)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 3)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 4)? 32'h1 : 
                                                   (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_inc_act_laddr_small = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_inc_act_laddr_large = (conv2d_25_control_param_index == 0)? 32'h3 : 
                                                (conv2d_25_control_param_index == 1)? 32'h10 : 
                                                (conv2d_25_control_param_index == 2)? 32'h20 : 
                                                (conv2d_25_control_param_index == 3)? 32'h40 : 
                                                (conv2d_25_control_param_index == 4)? 32'h80 : 
                                                (conv2d_25_control_param_index == 5)? 32'h100 : 32'h200;
  assign cparam_conv2d_25_inc_out_laddr_col = (conv2d_25_control_param_index == 0)? 32'h10 : 
                                              (conv2d_25_control_param_index == 1)? 32'h20 : 
                                              (conv2d_25_control_param_index == 2)? 32'h40 : 
                                              (conv2d_25_control_param_index == 3)? 32'h80 : 
                                              (conv2d_25_control_param_index == 4)? 32'h100 : 
                                              (conv2d_25_control_param_index == 5)? 32'h200 : 32'h400;
  assign cparam_conv2d_25_stream_act_local_small_offset = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                          (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                          (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                          (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                          (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                          (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_stream_act_local_large_offset = (conv2d_25_control_param_index == 0)? -32'sh3 : 
                                                          (conv2d_25_control_param_index == 1)? -32'sh10 : 
                                                          (conv2d_25_control_param_index == 2)? -32'sh20 : 
                                                          (conv2d_25_control_param_index == 3)? -32'sh40 : 
                                                          (conv2d_25_control_param_index == 4)? -32'sh80 : 
                                                          (conv2d_25_control_param_index == 5)? -32'sh100 : -32'sh200;
  assign cparam_conv2d_25_stream_act_local_small_flags_0 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_stream_act_local_small_flags_1 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_stream_act_local_small_flags_2 = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                                           (conv2d_25_control_param_index == 1)? 32'h1 : 
                                                           (conv2d_25_control_param_index == 2)? 32'h1 : 
                                                           (conv2d_25_control_param_index == 3)? 32'h1 : 
                                                           (conv2d_25_control_param_index == 4)? 32'h1 : 
                                                           (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_stream_act_local_large_flags_0 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_stream_act_local_large_flags_1 = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 1)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 2)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 3)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 4)? 32'h0 : 
                                                           (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  assign cparam_conv2d_25_stream_act_local_large_flags_2 = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                                           (conv2d_25_control_param_index == 1)? 32'h1 : 
                                                           (conv2d_25_control_param_index == 2)? 32'h1 : 
                                                           (conv2d_25_control_param_index == 3)? 32'h1 : 
                                                           (conv2d_25_control_param_index == 4)? 32'h1 : 
                                                           (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_inc_sync_out = (conv2d_25_control_param_index == 0)? 32'h1 : 
                                         (conv2d_25_control_param_index == 1)? 32'h1 : 
                                         (conv2d_25_control_param_index == 2)? 32'h1 : 
                                         (conv2d_25_control_param_index == 3)? 32'h1 : 
                                         (conv2d_25_control_param_index == 4)? 32'h1 : 
                                         (conv2d_25_control_param_index == 5)? 32'h1 : 32'h1;
  assign cparam_conv2d_25_inc_sync_out_res = (conv2d_25_control_param_index == 0)? 32'h0 : 
                                             (conv2d_25_control_param_index == 1)? 32'h0 : 
                                             (conv2d_25_control_param_index == 2)? 32'h0 : 
                                             (conv2d_25_control_param_index == 3)? 32'h0 : 
                                             (conv2d_25_control_param_index == 4)? 32'h0 : 
                                             (conv2d_25_control_param_index == 5)? 32'h0 : 32'h0;
  wire [9-1:0] cparam_max_pool_serial_27_act_num_col;
  wire [9-1:0] cparam_max_pool_serial_27_act_num_row;
  wire [2-1:0] cparam_max_pool_serial_27_stride_col;
  wire [2-1:0] cparam_max_pool_serial_27_stride_row;
  wire [8-1:0] cparam_max_pool_serial_27_out_num_col;
  wire [8-1:0] cparam_max_pool_serial_27_out_num_row;
  wire [1-1:0] cparam_max_pool_serial_27_pad_col_left;
  wire [1-1:0] cparam_max_pool_serial_27_pad_row_top;
  wire [9-1:0] cparam_max_pool_serial_27_max_col_count;
  wire [9-1:0] cparam_max_pool_serial_27_max_row_count;
  wire [1-1:0] cparam_max_pool_serial_27_max_bat_count;
  wire signed [32-1:0] cparam_max_pool_serial_27_act_offset_values_0;
  wire signed [32-1:0] cparam_max_pool_serial_27_act_offset_values_1;
  wire [16-1:0] cparam_max_pool_serial_27_act_row_step;
  wire [24-1:0] cparam_max_pool_serial_27_act_bat_step;
  wire [13-1:0] cparam_max_pool_serial_27_act_read_size;
  wire [9-1:0] cparam_max_pool_serial_27_act_read_block;
  wire [14-1:0] cparam_max_pool_serial_27_out_row_step;
  wire [22-1:0] cparam_max_pool_serial_27_out_bat_step;
  wire [12-1:0] cparam_max_pool_serial_27_out_write_size;
  wire [9-1:0] cparam_max_pool_serial_27_stream_size;
  wire [1-1:0] cparam_max_pool_serial_27_col_select_initval;
  wire [1-1:0] cparam_max_pool_serial_27_stride_col_mod_ksize;
  wire [2-1:0] cparam_max_pool_serial_27_ksize_col_minus_stride_col_mod;
  wire [1-1:0] cparam_max_pool_serial_27_local_pad_offset;
  wire [10-1:0] cparam_max_pool_serial_27_inc_act_laddr;
  wire [9-1:0] cparam_max_pool_serial_27_inc_out_laddr;
  reg [3-1:0] max_pool_serial_27_control_param_index;
  assign cparam_max_pool_serial_27_act_num_col = (max_pool_serial_27_control_param_index == 0)? 32'h1a0 : 
                                                 (max_pool_serial_27_control_param_index == 1)? 32'hd0 : 
                                                 (max_pool_serial_27_control_param_index == 2)? 32'h68 : 
                                                 (max_pool_serial_27_control_param_index == 3)? 32'h34 : 32'h1a;
  assign cparam_max_pool_serial_27_act_num_row = (max_pool_serial_27_control_param_index == 0)? 32'h1a0 : 
                                                 (max_pool_serial_27_control_param_index == 1)? 32'hd0 : 
                                                 (max_pool_serial_27_control_param_index == 2)? 32'h68 : 
                                                 (max_pool_serial_27_control_param_index == 3)? 32'h34 : 32'h1a;
  assign cparam_max_pool_serial_27_stride_col = (max_pool_serial_27_control_param_index == 0)? 32'h2 : 
                                                (max_pool_serial_27_control_param_index == 1)? 32'h2 : 
                                                (max_pool_serial_27_control_param_index == 2)? 32'h2 : 
                                                (max_pool_serial_27_control_param_index == 3)? 32'h2 : 32'h2;
  assign cparam_max_pool_serial_27_stride_row = (max_pool_serial_27_control_param_index == 0)? 32'h2 : 
                                                (max_pool_serial_27_control_param_index == 1)? 32'h2 : 
                                                (max_pool_serial_27_control_param_index == 2)? 32'h2 : 
                                                (max_pool_serial_27_control_param_index == 3)? 32'h2 : 32'h2;
  assign cparam_max_pool_serial_27_out_num_col = (max_pool_serial_27_control_param_index == 0)? 32'hd0 : 
                                                 (max_pool_serial_27_control_param_index == 1)? 32'h68 : 
                                                 (max_pool_serial_27_control_param_index == 2)? 32'h34 : 
                                                 (max_pool_serial_27_control_param_index == 3)? 32'h1a : 32'hd;
  assign cparam_max_pool_serial_27_out_num_row = (max_pool_serial_27_control_param_index == 0)? 32'hd0 : 
                                                 (max_pool_serial_27_control_param_index == 1)? 32'h68 : 
                                                 (max_pool_serial_27_control_param_index == 2)? 32'h34 : 
                                                 (max_pool_serial_27_control_param_index == 3)? 32'h1a : 32'hd;
  assign cparam_max_pool_serial_27_pad_col_left = (max_pool_serial_27_control_param_index == 0)? 32'h0 : 
                                                  (max_pool_serial_27_control_param_index == 1)? 32'h0 : 
                                                  (max_pool_serial_27_control_param_index == 2)? 32'h0 : 
                                                  (max_pool_serial_27_control_param_index == 3)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_27_pad_row_top = (max_pool_serial_27_control_param_index == 0)? 32'h0 : 
                                                 (max_pool_serial_27_control_param_index == 1)? 32'h0 : 
                                                 (max_pool_serial_27_control_param_index == 2)? 32'h0 : 
                                                 (max_pool_serial_27_control_param_index == 3)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_27_max_col_count = (max_pool_serial_27_control_param_index == 0)? 32'h19d : 
                                                   (max_pool_serial_27_control_param_index == 1)? 32'hcd : 
                                                   (max_pool_serial_27_control_param_index == 2)? 32'h65 : 
                                                   (max_pool_serial_27_control_param_index == 3)? 32'h31 : 32'h17;
  assign cparam_max_pool_serial_27_max_row_count = (max_pool_serial_27_control_param_index == 0)? 32'h19d : 
                                                   (max_pool_serial_27_control_param_index == 1)? 32'hcd : 
                                                   (max_pool_serial_27_control_param_index == 2)? 32'h65 : 
                                                   (max_pool_serial_27_control_param_index == 3)? 32'h31 : 32'h17;
  assign cparam_max_pool_serial_27_max_bat_count = (max_pool_serial_27_control_param_index == 0)? 32'h0 : 
                                                   (max_pool_serial_27_control_param_index == 1)? 32'h0 : 
                                                   (max_pool_serial_27_control_param_index == 2)? 32'h0 : 
                                                   (max_pool_serial_27_control_param_index == 3)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_27_act_offset_values_0 = (max_pool_serial_27_control_param_index == 0)? 32'h0 : 
                                                         (max_pool_serial_27_control_param_index == 1)? 32'h0 : 
                                                         (max_pool_serial_27_control_param_index == 2)? 32'h0 : 
                                                         (max_pool_serial_27_control_param_index == 3)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_27_act_offset_values_1 = (max_pool_serial_27_control_param_index == 0)? 32'h6800 : 
                                                         (max_pool_serial_27_control_param_index == 1)? 32'h6800 : 
                                                         (max_pool_serial_27_control_param_index == 2)? 32'h6800 : 
                                                         (max_pool_serial_27_control_param_index == 3)? 32'h6800 : 32'h6800;
  assign cparam_max_pool_serial_27_act_row_step = (max_pool_serial_27_control_param_index == 0)? 32'hd000 : 
                                                  (max_pool_serial_27_control_param_index == 1)? 32'hd000 : 
                                                  (max_pool_serial_27_control_param_index == 2)? 32'hd000 : 
                                                  (max_pool_serial_27_control_param_index == 3)? 32'hd000 : 32'hd000;
  assign cparam_max_pool_serial_27_act_bat_step = (max_pool_serial_27_control_param_index == 0)? 32'ha90000 : 
                                                  (max_pool_serial_27_control_param_index == 1)? 32'h548000 : 
                                                  (max_pool_serial_27_control_param_index == 2)? 32'h2a4000 : 
                                                  (max_pool_serial_27_control_param_index == 3)? 32'h152000 : 32'ha9000;
  assign cparam_max_pool_serial_27_act_read_size = (max_pool_serial_27_control_param_index == 0)? 32'h1a00 : 
                                                   (max_pool_serial_27_control_param_index == 1)? 32'h1a00 : 
                                                   (max_pool_serial_27_control_param_index == 2)? 32'h1a00 : 
                                                   (max_pool_serial_27_control_param_index == 3)? 32'h1a00 : 32'h1a00;
  assign cparam_max_pool_serial_27_act_read_block = (max_pool_serial_27_control_param_index == 0)? 32'h10 : 
                                                    (max_pool_serial_27_control_param_index == 1)? 32'h20 : 
                                                    (max_pool_serial_27_control_param_index == 2)? 32'h40 : 
                                                    (max_pool_serial_27_control_param_index == 3)? 32'h80 : 32'h100;
  assign cparam_max_pool_serial_27_out_row_step = (max_pool_serial_27_control_param_index == 0)? 32'h3400 : 
                                                  (max_pool_serial_27_control_param_index == 1)? 32'h3400 : 
                                                  (max_pool_serial_27_control_param_index == 2)? 32'h3400 : 
                                                  (max_pool_serial_27_control_param_index == 3)? 32'h3400 : 32'h3400;
  assign cparam_max_pool_serial_27_out_bat_step = (max_pool_serial_27_control_param_index == 0)? 32'h2a4000 : 
                                                  (max_pool_serial_27_control_param_index == 1)? 32'h152000 : 
                                                  (max_pool_serial_27_control_param_index == 2)? 32'ha9000 : 
                                                  (max_pool_serial_27_control_param_index == 3)? 32'h54800 : 32'h2a400;
  assign cparam_max_pool_serial_27_out_write_size = (max_pool_serial_27_control_param_index == 0)? 32'hd00 : 
                                                    (max_pool_serial_27_control_param_index == 1)? 32'hd00 : 
                                                    (max_pool_serial_27_control_param_index == 2)? 32'hd00 : 
                                                    (max_pool_serial_27_control_param_index == 3)? 32'hd00 : 32'hd00;
  assign cparam_max_pool_serial_27_stream_size = (max_pool_serial_27_control_param_index == 0)? 32'h10 : 
                                                 (max_pool_serial_27_control_param_index == 1)? 32'h20 : 
                                                 (max_pool_serial_27_control_param_index == 2)? 32'h40 : 
                                                 (max_pool_serial_27_control_param_index == 3)? 32'h80 : 32'h100;
  assign cparam_max_pool_serial_27_col_select_initval = (max_pool_serial_27_control_param_index == 0)? 32'h0 : 
                                                        (max_pool_serial_27_control_param_index == 1)? 32'h0 : 
                                                        (max_pool_serial_27_control_param_index == 2)? 32'h0 : 
                                                        (max_pool_serial_27_control_param_index == 3)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_27_stride_col_mod_ksize = (max_pool_serial_27_control_param_index == 0)? 32'h0 : 
                                                          (max_pool_serial_27_control_param_index == 1)? 32'h0 : 
                                                          (max_pool_serial_27_control_param_index == 2)? 32'h0 : 
                                                          (max_pool_serial_27_control_param_index == 3)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_27_ksize_col_minus_stride_col_mod = (max_pool_serial_27_control_param_index == 0)? 32'h2 : 
                                                                    (max_pool_serial_27_control_param_index == 1)? 32'h2 : 
                                                                    (max_pool_serial_27_control_param_index == 2)? 32'h2 : 
                                                                    (max_pool_serial_27_control_param_index == 3)? 32'h2 : 32'h2;
  assign cparam_max_pool_serial_27_local_pad_offset = (max_pool_serial_27_control_param_index == 0)? 32'h0 : 
                                                      (max_pool_serial_27_control_param_index == 1)? 32'h0 : 
                                                      (max_pool_serial_27_control_param_index == 2)? 32'h0 : 
                                                      (max_pool_serial_27_control_param_index == 3)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_27_inc_act_laddr = (max_pool_serial_27_control_param_index == 0)? 32'h20 : 
                                                   (max_pool_serial_27_control_param_index == 1)? 32'h40 : 
                                                   (max_pool_serial_27_control_param_index == 2)? 32'h80 : 
                                                   (max_pool_serial_27_control_param_index == 3)? 32'h100 : 32'h200;
  assign cparam_max_pool_serial_27_inc_out_laddr = (max_pool_serial_27_control_param_index == 0)? 32'h10 : 
                                                   (max_pool_serial_27_control_param_index == 1)? 32'h20 : 
                                                   (max_pool_serial_27_control_param_index == 2)? 32'h40 : 
                                                   (max_pool_serial_27_control_param_index == 3)? 32'h80 : 32'h100;
  wire [4-1:0] cparam_max_pool_47_act_num_col;
  wire [4-1:0] cparam_max_pool_47_act_num_row;
  wire [1-1:0] cparam_max_pool_47_stride_col;
  wire [1-1:0] cparam_max_pool_47_stride_row;
  wire [4-1:0] cparam_max_pool_47_out_num_col;
  wire [4-1:0] cparam_max_pool_47_out_num_row;
  wire [1-1:0] cparam_max_pool_47_pad_col_left;
  wire [1-1:0] cparam_max_pool_47_pad_row_top;
  wire [4-1:0] cparam_max_pool_47_max_col_count;
  wire [4-1:0] cparam_max_pool_47_max_row_count;
  wire [1-1:0] cparam_max_pool_47_max_bat_count;
  wire [1-1:0] cparam_max_pool_47_dma_flag_conds_0;
  wire [1-1:0] cparam_max_pool_47_dma_flag_conds_1;
  wire signed [32-1:0] cparam_max_pool_47_act_offset_values_0;
  wire signed [32-1:0] cparam_max_pool_47_act_offset_values_1;
  wire [15-1:0] cparam_max_pool_47_act_row_step;
  wire [19-1:0] cparam_max_pool_47_act_bat_step;
  wire [13-1:0] cparam_max_pool_47_act_read_size;
  wire [10-1:0] cparam_max_pool_47_act_read_block;
  wire [15-1:0] cparam_max_pool_47_out_row_step;
  wire [19-1:0] cparam_max_pool_47_out_bat_step;
  wire [13-1:0] cparam_max_pool_47_out_write_size;
  wire [10-1:0] cparam_max_pool_47_stream_size;
  wire [1-1:0] cparam_max_pool_47_col_select_initval;
  wire [1-1:0] cparam_max_pool_47_stride_col_mod_ksize;
  wire [1-1:0] cparam_max_pool_47_ksize_col_minus_stride_col_mod;
  wire [1-1:0] cparam_max_pool_47_inc_act_laddr_conds_0;
  wire [1-1:0] cparam_max_pool_47_inc_act_laddr_conds_1;
  wire [1-1:0] cparam_max_pool_47_inc_act_laddr_conds_2;
  wire [1-1:0] cparam_max_pool_47_inc_act_laddr_conds_3;
  wire [1-1:0] cparam_max_pool_47_inc_act_laddr_conds_4;
  wire [1-1:0] cparam_max_pool_47_inc_act_laddr_conds_5;
  wire [1-1:0] cparam_max_pool_47_inc_act_laddr_conds_6;
  wire [1-1:0] cparam_max_pool_47_inc_act_laddr_conds_7;
  wire [1-1:0] cparam_max_pool_47_inc_act_laddr_small;
  wire [10-1:0] cparam_max_pool_47_inc_act_laddr_large;
  wire [10-1:0] cparam_max_pool_47_inc_out_laddr;
  wire [1-1:0] cparam_max_pool_47_stream_act_local_small_offset;
  wire [1-1:0] cparam_max_pool_47_stream_act_local_large_offset;
  wire [1-1:0] cparam_max_pool_47_stream_act_local_small_flags_0;
  wire [1-1:0] cparam_max_pool_47_stream_act_local_small_flags_1;
  wire [1-1:0] cparam_max_pool_47_stream_act_local_large_flags_0;
  wire [1-1:0] cparam_max_pool_47_stream_act_local_large_flags_1;
  assign cparam_max_pool_47_act_num_col = 13;
  assign cparam_max_pool_47_act_num_row = 13;
  assign cparam_max_pool_47_stride_col = 1;
  assign cparam_max_pool_47_stride_row = 1;
  assign cparam_max_pool_47_out_num_col = 12;
  assign cparam_max_pool_47_out_num_row = 12;
  assign cparam_max_pool_47_pad_col_left = 0;
  assign cparam_max_pool_47_pad_row_top = 0;
  assign cparam_max_pool_47_max_col_count = 11;
  assign cparam_max_pool_47_max_row_count = 11;
  assign cparam_max_pool_47_max_bat_count = 0;
  assign cparam_max_pool_47_dma_flag_conds_0 = 1;
  assign cparam_max_pool_47_dma_flag_conds_1 = 0;
  assign cparam_max_pool_47_act_offset_values_0 = 0;
  assign cparam_max_pool_47_act_offset_values_1 = 26624;
  assign cparam_max_pool_47_act_row_step = 26624;
  assign cparam_max_pool_47_act_bat_step = 346112;
  assign cparam_max_pool_47_act_read_size = 6656;
  assign cparam_max_pool_47_act_read_block = 512;
  assign cparam_max_pool_47_out_row_step = 24576;
  assign cparam_max_pool_47_out_bat_step = 294912;
  assign cparam_max_pool_47_out_write_size = 6144;
  assign cparam_max_pool_47_stream_size = 512;
  assign cparam_max_pool_47_col_select_initval = 0;
  assign cparam_max_pool_47_stride_col_mod_ksize = 1;
  assign cparam_max_pool_47_ksize_col_minus_stride_col_mod = 1;
  assign cparam_max_pool_47_inc_act_laddr_conds_0 = 1;
  assign cparam_max_pool_47_inc_act_laddr_conds_1 = 0;
  assign cparam_max_pool_47_inc_act_laddr_conds_2 = 0;
  assign cparam_max_pool_47_inc_act_laddr_conds_3 = 1;
  assign cparam_max_pool_47_inc_act_laddr_conds_4 = 1;
  assign cparam_max_pool_47_inc_act_laddr_conds_5 = 0;
  assign cparam_max_pool_47_inc_act_laddr_conds_6 = 0;
  assign cparam_max_pool_47_inc_act_laddr_conds_7 = 1;
  assign cparam_max_pool_47_inc_act_laddr_small = 0;
  assign cparam_max_pool_47_inc_act_laddr_large = 512;
  assign cparam_max_pool_47_inc_out_laddr = 512;
  assign cparam_max_pool_47_stream_act_local_small_offset = 0;
  assign cparam_max_pool_47_stream_act_local_large_offset = 0;
  assign cparam_max_pool_47_stream_act_local_small_flags_0 = 0;
  assign cparam_max_pool_47_stream_act_local_small_flags_1 = 0;
  assign cparam_max_pool_47_stream_act_local_large_flags_0 = 0;
  assign cparam_max_pool_47_stream_act_local_large_flags_1 = 0;
  reg __max_0_stream_ivalid;
  wire __max_0_stream_oready;
  wire __max_0_stream_internal_oready;
  assign __max_0_stream_internal_oready = 1;
  reg [32-1:0] __max_0_fsm;
  localparam __max_0_fsm_init = 0;
  wire __max_0_run_flag;
  assign __max_0_run_flag = 0;
  reg __max_0_source_start;
  wire __max_0_source_stop;
  reg __max_0_source_busy;
  wire __max_0_sink_start;
  wire __max_0_sink_stop;
  wire __max_0_sink_busy;
  wire __max_0_busy;
  reg __max_0_busy_reg;
  wire __max_0_is_root;
  reg __max_0_var0_idle;
  reg [33-1:0] __max_0_var0_source_count;
  reg [5-1:0] __max_0_var0_source_mode;
  reg [16-1:0] __max_0_var0_source_generator_id;
  reg [32-1:0] __max_0_var0_source_offset;
  reg [33-1:0] __max_0_var0_source_size;
  reg [32-1:0] __max_0_var0_source_stride;
  reg [32-1:0] __max_0_var0_source_offset_buf;
  reg [33-1:0] __max_0_var0_source_size_buf;
  reg [32-1:0] __max_0_var0_source_stride_buf;
  reg [8-1:0] __max_0_var0_source_sel;
  reg [32-1:0] __max_0_var0_source_ram_raddr;
  reg __max_0_var0_source_ram_renable;
  wire [32-1:0] __max_0_var0_source_ram_rdata;
  reg __max_0_var0_source_fifo_deq;
  wire [32-1:0] __max_0_var0_source_fifo_rdata;
  reg [32-1:0] __max_0_var0_source_empty_data;
  reg __max_0_var1_idle;
  reg [33-1:0] __max_0_var1_source_count;
  reg [5-1:0] __max_0_var1_source_mode;
  reg [16-1:0] __max_0_var1_source_generator_id;
  reg [32-1:0] __max_0_var1_source_offset;
  reg [33-1:0] __max_0_var1_source_size;
  reg [32-1:0] __max_0_var1_source_stride;
  reg [32-1:0] __max_0_var1_source_offset_buf;
  reg [33-1:0] __max_0_var1_source_size_buf;
  reg [32-1:0] __max_0_var1_source_stride_buf;
  reg [8-1:0] __max_0_var1_source_sel;
  reg [32-1:0] __max_0_var1_source_ram_raddr;
  reg __max_0_var1_source_ram_renable;
  wire [32-1:0] __max_0_var1_source_ram_rdata;
  reg __max_0_var1_source_fifo_deq;
  wire [32-1:0] __max_0_var1_source_fifo_rdata;
  reg [32-1:0] __max_0_var1_source_empty_data;
  reg __max_0_var2_idle;
  reg [33-1:0] __max_0_var2_source_count;
  reg [5-1:0] __max_0_var2_source_mode;
  reg [16-1:0] __max_0_var2_source_generator_id;
  reg [32-1:0] __max_0_var2_source_offset;
  reg [33-1:0] __max_0_var2_source_size;
  reg [32-1:0] __max_0_var2_source_stride;
  reg [32-1:0] __max_0_var2_source_offset_buf;
  reg [33-1:0] __max_0_var2_source_size_buf;
  reg [32-1:0] __max_0_var2_source_stride_buf;
  reg [8-1:0] __max_0_var2_source_sel;
  reg [32-1:0] __max_0_var2_source_ram_raddr;
  reg __max_0_var2_source_ram_renable;
  wire [32-1:0] __max_0_var2_source_ram_rdata;
  reg __max_0_var2_source_fifo_deq;
  wire [32-1:0] __max_0_var2_source_fifo_rdata;
  reg [32-1:0] __max_0_var2_source_empty_data;
  reg __max_0_var3_idle;
  reg [33-1:0] __max_0_var3_source_count;
  reg [5-1:0] __max_0_var3_source_mode;
  reg [16-1:0] __max_0_var3_source_generator_id;
  reg [32-1:0] __max_0_var3_source_offset;
  reg [33-1:0] __max_0_var3_source_size;
  reg [32-1:0] __max_0_var3_source_stride;
  reg [32-1:0] __max_0_var3_source_offset_buf;
  reg [33-1:0] __max_0_var3_source_size_buf;
  reg [32-1:0] __max_0_var3_source_stride_buf;
  reg [8-1:0] __max_0_var3_source_sel;
  reg [32-1:0] __max_0_var3_source_ram_raddr;
  reg __max_0_var3_source_ram_renable;
  wire [32-1:0] __max_0_var3_source_ram_rdata;
  reg __max_0_var3_source_fifo_deq;
  wire [32-1:0] __max_0_var3_source_fifo_rdata;
  reg [32-1:0] __max_0_var3_source_empty_data;
  reg [33-1:0] __max_0_val_sink_count;
  reg [5-1:0] __max_0_val_sink_mode;
  reg [16-1:0] __max_0_val_sink_generator_id;
  reg [32-1:0] __max_0_val_sink_offset;
  reg [33-1:0] __max_0_val_sink_size;
  reg [32-1:0] __max_0_val_sink_stride;
  reg [32-1:0] __max_0_val_sink_offset_buf;
  reg [33-1:0] __max_0_val_sink_size_buf;
  reg [32-1:0] __max_0_val_sink_stride_buf;
  reg [8-1:0] __max_0_val_sink_sel;
  reg [32-1:0] __max_0_val_sink_waddr;
  reg __max_0_val_sink_wenable;
  reg [32-1:0] __max_0_val_sink_wdata;
  reg __max_0_val_sink_fifo_enq;
  reg [32-1:0] __max_0_val_sink_fifo_wdata;
  reg [32-1:0] __max_0_val_sink_immediate;
  reg _acc_1_stream_ivalid;
  wire _acc_1_stream_oready;
  wire _acc_1_stream_internal_oready;
  assign _acc_1_stream_internal_oready = 1;
  reg [32-1:0] _acc_1_fsm;
  localparam _acc_1_fsm_init = 0;
  wire _acc_1_run_flag;
  assign _acc_1_run_flag = 0;
  reg _acc_1_source_start;
  wire _acc_1_source_stop;
  reg _acc_1_source_busy;
  wire _acc_1_sink_start;
  wire _acc_1_sink_stop;
  wire _acc_1_sink_busy;
  wire _acc_1_busy;
  reg _acc_1_busy_reg;
  wire _acc_1_is_root;
  reg _acc_1_x_idle;
  reg [33-1:0] _acc_1_x_source_count;
  reg [5-1:0] _acc_1_x_source_mode;
  reg [16-1:0] _acc_1_x_source_generator_id;
  reg [32-1:0] _acc_1_x_source_offset;
  reg [33-1:0] _acc_1_x_source_size;
  reg [32-1:0] _acc_1_x_source_stride;
  reg [32-1:0] _acc_1_x_source_offset_buf;
  reg [33-1:0] _acc_1_x_source_size_buf;
  reg [32-1:0] _acc_1_x_source_stride_buf;
  reg [8-1:0] _acc_1_x_source_sel;
  reg [32-1:0] _acc_1_x_source_ram_raddr;
  reg _acc_1_x_source_ram_renable;
  wire [128-1:0] _acc_1_x_source_ram_rdata;
  reg _acc_1_x_source_fifo_deq;
  wire [128-1:0] _acc_1_x_source_fifo_rdata;
  reg [128-1:0] _acc_1_x_source_empty_data;
  reg _acc_1_rshift_idle;
  reg [33-1:0] _acc_1_rshift_source_count;
  reg [5-1:0] _acc_1_rshift_source_mode;
  reg [16-1:0] _acc_1_rshift_source_generator_id;
  reg [32-1:0] _acc_1_rshift_source_offset;
  reg [33-1:0] _acc_1_rshift_source_size;
  reg [32-1:0] _acc_1_rshift_source_stride;
  reg [32-1:0] _acc_1_rshift_source_offset_buf;
  reg [33-1:0] _acc_1_rshift_source_size_buf;
  reg [32-1:0] _acc_1_rshift_source_stride_buf;
  reg [8-1:0] _acc_1_rshift_source_sel;
  reg [32-1:0] _acc_1_rshift_source_ram_raddr;
  reg _acc_1_rshift_source_ram_renable;
  wire [32-1:0] _acc_1_rshift_source_ram_rdata;
  reg _acc_1_rshift_source_fifo_deq;
  wire [32-1:0] _acc_1_rshift_source_fifo_rdata;
  reg [32-1:0] _acc_1_rshift_source_empty_data;
  reg [32-1:0] _acc_1_size_next_parameter_data;
  reg [33-1:0] _acc_1_sum_sink_count;
  reg [5-1:0] _acc_1_sum_sink_mode;
  reg [16-1:0] _acc_1_sum_sink_generator_id;
  reg [32-1:0] _acc_1_sum_sink_offset;
  reg [33-1:0] _acc_1_sum_sink_size;
  reg [32-1:0] _acc_1_sum_sink_stride;
  reg [32-1:0] _acc_1_sum_sink_offset_buf;
  reg [33-1:0] _acc_1_sum_sink_size_buf;
  reg [32-1:0] _acc_1_sum_sink_stride_buf;
  reg [8-1:0] _acc_1_sum_sink_sel;
  reg [32-1:0] _acc_1_sum_sink_waddr;
  reg _acc_1_sum_sink_wenable;
  reg [128-1:0] _acc_1_sum_sink_wdata;
  reg _acc_1_sum_sink_fifo_enq;
  reg [128-1:0] _acc_1_sum_sink_fifo_wdata;
  reg [128-1:0] _acc_1_sum_sink_immediate;
  reg [33-1:0] _acc_1_valid_sink_count;
  reg [5-1:0] _acc_1_valid_sink_mode;
  reg [16-1:0] _acc_1_valid_sink_generator_id;
  reg [32-1:0] _acc_1_valid_sink_offset;
  reg [33-1:0] _acc_1_valid_sink_size;
  reg [32-1:0] _acc_1_valid_sink_stride;
  reg [32-1:0] _acc_1_valid_sink_offset_buf;
  reg [33-1:0] _acc_1_valid_sink_size_buf;
  reg [32-1:0] _acc_1_valid_sink_stride_buf;
  reg [8-1:0] _acc_1_valid_sink_sel;
  reg [32-1:0] _acc_1_valid_sink_waddr;
  reg _acc_1_valid_sink_wenable;
  reg [1-1:0] _acc_1_valid_sink_wdata;
  reg _acc_1_valid_sink_fifo_enq;
  reg [1-1:0] _acc_1_valid_sink_fifo_wdata;
  reg [1-1:0] _acc_1_valid_sink_immediate;
  reg _add_tree_2_stream_ivalid;
  wire _add_tree_2_stream_oready;
  wire _add_tree_2_stream_internal_oready;
  assign _add_tree_2_stream_internal_oready = 1;
  reg [32-1:0] _add_tree_2_fsm;
  localparam _add_tree_2_fsm_init = 0;
  wire _add_tree_2_run_flag;
  assign _add_tree_2_run_flag = 0;
  reg _add_tree_2_source_start;
  wire _add_tree_2_source_stop;
  reg _add_tree_2_source_busy;
  wire _add_tree_2_sink_start;
  wire _add_tree_2_sink_stop;
  wire _add_tree_2_sink_busy;
  wire _add_tree_2_busy;
  reg _add_tree_2_busy_reg;
  wire _add_tree_2_is_root;
  reg _add_tree_2_var0_idle;
  reg [33-1:0] _add_tree_2_var0_source_count;
  reg [5-1:0] _add_tree_2_var0_source_mode;
  reg [16-1:0] _add_tree_2_var0_source_generator_id;
  reg [32-1:0] _add_tree_2_var0_source_offset;
  reg [33-1:0] _add_tree_2_var0_source_size;
  reg [32-1:0] _add_tree_2_var0_source_stride;
  reg [32-1:0] _add_tree_2_var0_source_offset_buf;
  reg [33-1:0] _add_tree_2_var0_source_size_buf;
  reg [32-1:0] _add_tree_2_var0_source_stride_buf;
  reg [8-1:0] _add_tree_2_var0_source_sel;
  reg [32-1:0] _add_tree_2_var0_source_ram_raddr;
  reg _add_tree_2_var0_source_ram_renable;
  wire [128-1:0] _add_tree_2_var0_source_ram_rdata;
  reg _add_tree_2_var0_source_fifo_deq;
  wire [128-1:0] _add_tree_2_var0_source_fifo_rdata;
  reg [128-1:0] _add_tree_2_var0_source_empty_data;
  reg _add_tree_2_var1_idle;
  reg [33-1:0] _add_tree_2_var1_source_count;
  reg [5-1:0] _add_tree_2_var1_source_mode;
  reg [16-1:0] _add_tree_2_var1_source_generator_id;
  reg [32-1:0] _add_tree_2_var1_source_offset;
  reg [33-1:0] _add_tree_2_var1_source_size;
  reg [32-1:0] _add_tree_2_var1_source_stride;
  reg [32-1:0] _add_tree_2_var1_source_offset_buf;
  reg [33-1:0] _add_tree_2_var1_source_size_buf;
  reg [32-1:0] _add_tree_2_var1_source_stride_buf;
  reg [8-1:0] _add_tree_2_var1_source_sel;
  reg [32-1:0] _add_tree_2_var1_source_ram_raddr;
  reg _add_tree_2_var1_source_ram_renable;
  wire [128-1:0] _add_tree_2_var1_source_ram_rdata;
  reg _add_tree_2_var1_source_fifo_deq;
  wire [128-1:0] _add_tree_2_var1_source_fifo_rdata;
  reg [128-1:0] _add_tree_2_var1_source_empty_data;
  reg _add_tree_2_var2_idle;
  reg [33-1:0] _add_tree_2_var2_source_count;
  reg [5-1:0] _add_tree_2_var2_source_mode;
  reg [16-1:0] _add_tree_2_var2_source_generator_id;
  reg [32-1:0] _add_tree_2_var2_source_offset;
  reg [33-1:0] _add_tree_2_var2_source_size;
  reg [32-1:0] _add_tree_2_var2_source_stride;
  reg [32-1:0] _add_tree_2_var2_source_offset_buf;
  reg [33-1:0] _add_tree_2_var2_source_size_buf;
  reg [32-1:0] _add_tree_2_var2_source_stride_buf;
  reg [8-1:0] _add_tree_2_var2_source_sel;
  reg [32-1:0] _add_tree_2_var2_source_ram_raddr;
  reg _add_tree_2_var2_source_ram_renable;
  wire [128-1:0] _add_tree_2_var2_source_ram_rdata;
  reg _add_tree_2_var2_source_fifo_deq;
  wire [128-1:0] _add_tree_2_var2_source_fifo_rdata;
  reg [128-1:0] _add_tree_2_var2_source_empty_data;
  reg _add_tree_2_var3_idle;
  reg [33-1:0] _add_tree_2_var3_source_count;
  reg [5-1:0] _add_tree_2_var3_source_mode;
  reg [16-1:0] _add_tree_2_var3_source_generator_id;
  reg [32-1:0] _add_tree_2_var3_source_offset;
  reg [33-1:0] _add_tree_2_var3_source_size;
  reg [32-1:0] _add_tree_2_var3_source_stride;
  reg [32-1:0] _add_tree_2_var3_source_offset_buf;
  reg [33-1:0] _add_tree_2_var3_source_size_buf;
  reg [32-1:0] _add_tree_2_var3_source_stride_buf;
  reg [8-1:0] _add_tree_2_var3_source_sel;
  reg [32-1:0] _add_tree_2_var3_source_ram_raddr;
  reg _add_tree_2_var3_source_ram_renable;
  wire [128-1:0] _add_tree_2_var3_source_ram_rdata;
  reg _add_tree_2_var3_source_fifo_deq;
  wire [128-1:0] _add_tree_2_var3_source_fifo_rdata;
  reg [128-1:0] _add_tree_2_var3_source_empty_data;
  reg _add_tree_2_var4_idle;
  reg [33-1:0] _add_tree_2_var4_source_count;
  reg [5-1:0] _add_tree_2_var4_source_mode;
  reg [16-1:0] _add_tree_2_var4_source_generator_id;
  reg [32-1:0] _add_tree_2_var4_source_offset;
  reg [33-1:0] _add_tree_2_var4_source_size;
  reg [32-1:0] _add_tree_2_var4_source_stride;
  reg [32-1:0] _add_tree_2_var4_source_offset_buf;
  reg [33-1:0] _add_tree_2_var4_source_size_buf;
  reg [32-1:0] _add_tree_2_var4_source_stride_buf;
  reg [8-1:0] _add_tree_2_var4_source_sel;
  reg [32-1:0] _add_tree_2_var4_source_ram_raddr;
  reg _add_tree_2_var4_source_ram_renable;
  wire [128-1:0] _add_tree_2_var4_source_ram_rdata;
  reg _add_tree_2_var4_source_fifo_deq;
  wire [128-1:0] _add_tree_2_var4_source_fifo_rdata;
  reg [128-1:0] _add_tree_2_var4_source_empty_data;
  reg _add_tree_2_var5_idle;
  reg [33-1:0] _add_tree_2_var5_source_count;
  reg [5-1:0] _add_tree_2_var5_source_mode;
  reg [16-1:0] _add_tree_2_var5_source_generator_id;
  reg [32-1:0] _add_tree_2_var5_source_offset;
  reg [33-1:0] _add_tree_2_var5_source_size;
  reg [32-1:0] _add_tree_2_var5_source_stride;
  reg [32-1:0] _add_tree_2_var5_source_offset_buf;
  reg [33-1:0] _add_tree_2_var5_source_size_buf;
  reg [32-1:0] _add_tree_2_var5_source_stride_buf;
  reg [8-1:0] _add_tree_2_var5_source_sel;
  reg [32-1:0] _add_tree_2_var5_source_ram_raddr;
  reg _add_tree_2_var5_source_ram_renable;
  wire [128-1:0] _add_tree_2_var5_source_ram_rdata;
  reg _add_tree_2_var5_source_fifo_deq;
  wire [128-1:0] _add_tree_2_var5_source_fifo_rdata;
  reg [128-1:0] _add_tree_2_var5_source_empty_data;
  reg _add_tree_2_var6_idle;
  reg [33-1:0] _add_tree_2_var6_source_count;
  reg [5-1:0] _add_tree_2_var6_source_mode;
  reg [16-1:0] _add_tree_2_var6_source_generator_id;
  reg [32-1:0] _add_tree_2_var6_source_offset;
  reg [33-1:0] _add_tree_2_var6_source_size;
  reg [32-1:0] _add_tree_2_var6_source_stride;
  reg [32-1:0] _add_tree_2_var6_source_offset_buf;
  reg [33-1:0] _add_tree_2_var6_source_size_buf;
  reg [32-1:0] _add_tree_2_var6_source_stride_buf;
  reg [8-1:0] _add_tree_2_var6_source_sel;
  reg [32-1:0] _add_tree_2_var6_source_ram_raddr;
  reg _add_tree_2_var6_source_ram_renable;
  wire [128-1:0] _add_tree_2_var6_source_ram_rdata;
  reg _add_tree_2_var6_source_fifo_deq;
  wire [128-1:0] _add_tree_2_var6_source_fifo_rdata;
  reg [128-1:0] _add_tree_2_var6_source_empty_data;
  reg _add_tree_2_var7_idle;
  reg [33-1:0] _add_tree_2_var7_source_count;
  reg [5-1:0] _add_tree_2_var7_source_mode;
  reg [16-1:0] _add_tree_2_var7_source_generator_id;
  reg [32-1:0] _add_tree_2_var7_source_offset;
  reg [33-1:0] _add_tree_2_var7_source_size;
  reg [32-1:0] _add_tree_2_var7_source_stride;
  reg [32-1:0] _add_tree_2_var7_source_offset_buf;
  reg [33-1:0] _add_tree_2_var7_source_size_buf;
  reg [32-1:0] _add_tree_2_var7_source_stride_buf;
  reg [8-1:0] _add_tree_2_var7_source_sel;
  reg [32-1:0] _add_tree_2_var7_source_ram_raddr;
  reg _add_tree_2_var7_source_ram_renable;
  wire [128-1:0] _add_tree_2_var7_source_ram_rdata;
  reg _add_tree_2_var7_source_fifo_deq;
  wire [128-1:0] _add_tree_2_var7_source_fifo_rdata;
  reg [128-1:0] _add_tree_2_var7_source_empty_data;
  reg _add_tree_2_var8_idle;
  reg [33-1:0] _add_tree_2_var8_source_count;
  reg [5-1:0] _add_tree_2_var8_source_mode;
  reg [16-1:0] _add_tree_2_var8_source_generator_id;
  reg [32-1:0] _add_tree_2_var8_source_offset;
  reg [33-1:0] _add_tree_2_var8_source_size;
  reg [32-1:0] _add_tree_2_var8_source_stride;
  reg [32-1:0] _add_tree_2_var8_source_offset_buf;
  reg [33-1:0] _add_tree_2_var8_source_size_buf;
  reg [32-1:0] _add_tree_2_var8_source_stride_buf;
  reg [8-1:0] _add_tree_2_var8_source_sel;
  reg [32-1:0] _add_tree_2_var8_source_ram_raddr;
  reg _add_tree_2_var8_source_ram_renable;
  wire [128-1:0] _add_tree_2_var8_source_ram_rdata;
  reg _add_tree_2_var8_source_fifo_deq;
  wire [128-1:0] _add_tree_2_var8_source_fifo_rdata;
  reg [128-1:0] _add_tree_2_var8_source_empty_data;
  reg [33-1:0] _add_tree_2_sum_sink_count;
  reg [5-1:0] _add_tree_2_sum_sink_mode;
  reg [16-1:0] _add_tree_2_sum_sink_generator_id;
  reg [32-1:0] _add_tree_2_sum_sink_offset;
  reg [33-1:0] _add_tree_2_sum_sink_size;
  reg [32-1:0] _add_tree_2_sum_sink_stride;
  reg [32-1:0] _add_tree_2_sum_sink_offset_buf;
  reg [33-1:0] _add_tree_2_sum_sink_size_buf;
  reg [32-1:0] _add_tree_2_sum_sink_stride_buf;
  reg [8-1:0] _add_tree_2_sum_sink_sel;
  reg [32-1:0] _add_tree_2_sum_sink_waddr;
  reg _add_tree_2_sum_sink_wenable;
  reg [128-1:0] _add_tree_2_sum_sink_wdata;
  reg _add_tree_2_sum_sink_fifo_enq;
  reg [128-1:0] _add_tree_2_sum_sink_fifo_wdata;
  reg [128-1:0] _add_tree_2_sum_sink_immediate;
  reg _mul_rshift_round_clip_3_stream_ivalid;
  wire _mul_rshift_round_clip_3_stream_oready;
  wire _mul_rshift_round_clip_3_stream_internal_oready;
  assign _mul_rshift_round_clip_3_stream_internal_oready = 1;
  reg [32-1:0] _mul_rshift_round_clip_3_fsm;
  localparam _mul_rshift_round_clip_3_fsm_init = 0;
  wire _mul_rshift_round_clip_3_run_flag;
  assign _mul_rshift_round_clip_3_run_flag = 0;
  reg _mul_rshift_round_clip_3_source_start;
  wire _mul_rshift_round_clip_3_source_stop;
  reg _mul_rshift_round_clip_3_source_busy;
  wire _mul_rshift_round_clip_3_sink_start;
  wire _mul_rshift_round_clip_3_sink_stop;
  wire _mul_rshift_round_clip_3_sink_busy;
  wire _mul_rshift_round_clip_3_busy;
  reg _mul_rshift_round_clip_3_busy_reg;
  wire _mul_rshift_round_clip_3_is_root;
  reg _mul_rshift_round_clip_3_x_idle;
  reg [33-1:0] _mul_rshift_round_clip_3_x_source_count;
  reg [5-1:0] _mul_rshift_round_clip_3_x_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_3_x_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_3_x_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_3_x_source_size;
  reg [32-1:0] _mul_rshift_round_clip_3_x_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_3_x_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_3_x_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_3_x_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_3_x_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_3_x_source_ram_raddr;
  reg _mul_rshift_round_clip_3_x_source_ram_renable;
  wire [128-1:0] _mul_rshift_round_clip_3_x_source_ram_rdata;
  reg _mul_rshift_round_clip_3_x_source_fifo_deq;
  wire [128-1:0] _mul_rshift_round_clip_3_x_source_fifo_rdata;
  reg [128-1:0] _mul_rshift_round_clip_3_x_source_empty_data;
  reg _mul_rshift_round_clip_3_y_idle;
  reg [33-1:0] _mul_rshift_round_clip_3_y_source_count;
  reg [5-1:0] _mul_rshift_round_clip_3_y_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_3_y_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_3_y_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_3_y_source_size;
  reg [32-1:0] _mul_rshift_round_clip_3_y_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_3_y_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_3_y_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_3_y_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_3_y_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_3_y_source_ram_raddr;
  reg _mul_rshift_round_clip_3_y_source_ram_renable;
  wire [32-1:0] _mul_rshift_round_clip_3_y_source_ram_rdata;
  reg _mul_rshift_round_clip_3_y_source_fifo_deq;
  wire [32-1:0] _mul_rshift_round_clip_3_y_source_fifo_rdata;
  reg [32-1:0] _mul_rshift_round_clip_3_y_source_empty_data;
  reg _mul_rshift_round_clip_3_rshift_idle;
  reg [33-1:0] _mul_rshift_round_clip_3_rshift_source_count;
  reg [5-1:0] _mul_rshift_round_clip_3_rshift_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_3_rshift_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_3_rshift_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_3_rshift_source_size;
  reg [32-1:0] _mul_rshift_round_clip_3_rshift_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_3_rshift_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_3_rshift_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_3_rshift_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_3_rshift_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_3_rshift_source_ram_raddr;
  reg _mul_rshift_round_clip_3_rshift_source_ram_renable;
  wire [32-1:0] _mul_rshift_round_clip_3_rshift_source_ram_rdata;
  reg _mul_rshift_round_clip_3_rshift_source_fifo_deq;
  wire [32-1:0] _mul_rshift_round_clip_3_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_rshift_round_clip_3_rshift_source_empty_data;
  reg [33-1:0] _mul_rshift_round_clip_3_z_sink_count;
  reg [5-1:0] _mul_rshift_round_clip_3_z_sink_mode;
  reg [16-1:0] _mul_rshift_round_clip_3_z_sink_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_3_z_sink_offset;
  reg [33-1:0] _mul_rshift_round_clip_3_z_sink_size;
  reg [32-1:0] _mul_rshift_round_clip_3_z_sink_stride;
  reg [32-1:0] _mul_rshift_round_clip_3_z_sink_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_3_z_sink_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_3_z_sink_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_3_z_sink_sel;
  reg [32-1:0] _mul_rshift_round_clip_3_z_sink_waddr;
  reg _mul_rshift_round_clip_3_z_sink_wenable;
  reg [32-1:0] _mul_rshift_round_clip_3_z_sink_wdata;
  reg _mul_rshift_round_clip_3_z_sink_fifo_enq;
  reg [32-1:0] _mul_rshift_round_clip_3_z_sink_fifo_wdata;
  reg [32-1:0] _mul_rshift_round_clip_3_z_sink_immediate;
  reg _mul_4_stream_ivalid;
  wire _mul_4_stream_oready;
  wire _mul_4_stream_internal_oready;
  assign _mul_4_stream_internal_oready = 1;
  reg [32-1:0] _mul_4_fsm;
  localparam _mul_4_fsm_init = 0;
  wire _mul_4_run_flag;
  assign _mul_4_run_flag = 0;
  reg _mul_4_source_start;
  wire _mul_4_source_stop;
  reg _mul_4_source_busy;
  wire _mul_4_sink_start;
  wire _mul_4_sink_stop;
  wire _mul_4_sink_busy;
  wire _mul_4_busy;
  reg _mul_4_busy_reg;
  wire _mul_4_is_root;
  reg _mul_4_x_idle;
  reg [33-1:0] _mul_4_x_source_count;
  reg [5-1:0] _mul_4_x_source_mode;
  reg [16-1:0] _mul_4_x_source_generator_id;
  reg [32-1:0] _mul_4_x_source_offset;
  reg [33-1:0] _mul_4_x_source_size;
  reg [32-1:0] _mul_4_x_source_stride;
  reg [32-1:0] _mul_4_x_source_offset_buf;
  reg [33-1:0] _mul_4_x_source_size_buf;
  reg [32-1:0] _mul_4_x_source_stride_buf;
  reg [8-1:0] _mul_4_x_source_sel;
  reg [32-1:0] _mul_4_x_source_ram_raddr;
  reg _mul_4_x_source_ram_renable;
  wire [32-1:0] _mul_4_x_source_ram_rdata;
  reg _mul_4_x_source_fifo_deq;
  wire [32-1:0] _mul_4_x_source_fifo_rdata;
  reg [32-1:0] _mul_4_x_source_empty_data;
  reg _mul_4_y_idle;
  reg [33-1:0] _mul_4_y_source_count;
  reg [5-1:0] _mul_4_y_source_mode;
  reg [16-1:0] _mul_4_y_source_generator_id;
  reg [32-1:0] _mul_4_y_source_offset;
  reg [33-1:0] _mul_4_y_source_size;
  reg [32-1:0] _mul_4_y_source_stride;
  reg [32-1:0] _mul_4_y_source_offset_buf;
  reg [33-1:0] _mul_4_y_source_size_buf;
  reg [32-1:0] _mul_4_y_source_stride_buf;
  reg [8-1:0] _mul_4_y_source_sel;
  reg [32-1:0] _mul_4_y_source_ram_raddr;
  reg _mul_4_y_source_ram_renable;
  wire [32-1:0] _mul_4_y_source_ram_rdata;
  reg _mul_4_y_source_fifo_deq;
  wire [32-1:0] _mul_4_y_source_fifo_rdata;
  reg [32-1:0] _mul_4_y_source_empty_data;
  reg _mul_4_rshift_idle;
  reg [33-1:0] _mul_4_rshift_source_count;
  reg [5-1:0] _mul_4_rshift_source_mode;
  reg [16-1:0] _mul_4_rshift_source_generator_id;
  reg [32-1:0] _mul_4_rshift_source_offset;
  reg [33-1:0] _mul_4_rshift_source_size;
  reg [32-1:0] _mul_4_rshift_source_stride;
  reg [32-1:0] _mul_4_rshift_source_offset_buf;
  reg [33-1:0] _mul_4_rshift_source_size_buf;
  reg [32-1:0] _mul_4_rshift_source_stride_buf;
  reg [8-1:0] _mul_4_rshift_source_sel;
  reg [32-1:0] _mul_4_rshift_source_ram_raddr;
  reg _mul_4_rshift_source_ram_renable;
  wire [32-1:0] _mul_4_rshift_source_ram_rdata;
  reg _mul_4_rshift_source_fifo_deq;
  wire [32-1:0] _mul_4_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_4_rshift_source_empty_data;
  reg [33-1:0] _mul_4_z_sink_count;
  reg [5-1:0] _mul_4_z_sink_mode;
  reg [16-1:0] _mul_4_z_sink_generator_id;
  reg [32-1:0] _mul_4_z_sink_offset;
  reg [33-1:0] _mul_4_z_sink_size;
  reg [32-1:0] _mul_4_z_sink_stride;
  reg [32-1:0] _mul_4_z_sink_offset_buf;
  reg [33-1:0] _mul_4_z_sink_size_buf;
  reg [32-1:0] _mul_4_z_sink_stride_buf;
  reg [8-1:0] _mul_4_z_sink_sel;
  reg [32-1:0] _mul_4_z_sink_waddr;
  reg _mul_4_z_sink_wenable;
  reg [64-1:0] _mul_4_z_sink_wdata;
  reg _mul_4_z_sink_fifo_enq;
  reg [64-1:0] _mul_4_z_sink_fifo_wdata;
  reg [64-1:0] _mul_4_z_sink_immediate;
  reg _mul_5_stream_ivalid;
  wire _mul_5_stream_oready;
  wire _mul_5_stream_internal_oready;
  assign _mul_5_stream_internal_oready = 1;
  reg [32-1:0] _mul_5_fsm;
  localparam _mul_5_fsm_init = 0;
  wire _mul_5_run_flag;
  assign _mul_5_run_flag = 0;
  reg _mul_5_source_start;
  wire _mul_5_source_stop;
  reg _mul_5_source_busy;
  wire _mul_5_sink_start;
  wire _mul_5_sink_stop;
  wire _mul_5_sink_busy;
  wire _mul_5_busy;
  reg _mul_5_busy_reg;
  wire _mul_5_is_root;
  reg _mul_5_x_idle;
  reg [33-1:0] _mul_5_x_source_count;
  reg [5-1:0] _mul_5_x_source_mode;
  reg [16-1:0] _mul_5_x_source_generator_id;
  reg [32-1:0] _mul_5_x_source_offset;
  reg [33-1:0] _mul_5_x_source_size;
  reg [32-1:0] _mul_5_x_source_stride;
  reg [32-1:0] _mul_5_x_source_offset_buf;
  reg [33-1:0] _mul_5_x_source_size_buf;
  reg [32-1:0] _mul_5_x_source_stride_buf;
  reg [8-1:0] _mul_5_x_source_sel;
  reg [32-1:0] _mul_5_x_source_ram_raddr;
  reg _mul_5_x_source_ram_renable;
  wire [32-1:0] _mul_5_x_source_ram_rdata;
  reg _mul_5_x_source_fifo_deq;
  wire [32-1:0] _mul_5_x_source_fifo_rdata;
  reg [32-1:0] _mul_5_x_source_empty_data;
  reg _mul_5_y_idle;
  reg [33-1:0] _mul_5_y_source_count;
  reg [5-1:0] _mul_5_y_source_mode;
  reg [16-1:0] _mul_5_y_source_generator_id;
  reg [32-1:0] _mul_5_y_source_offset;
  reg [33-1:0] _mul_5_y_source_size;
  reg [32-1:0] _mul_5_y_source_stride;
  reg [32-1:0] _mul_5_y_source_offset_buf;
  reg [33-1:0] _mul_5_y_source_size_buf;
  reg [32-1:0] _mul_5_y_source_stride_buf;
  reg [8-1:0] _mul_5_y_source_sel;
  reg [32-1:0] _mul_5_y_source_ram_raddr;
  reg _mul_5_y_source_ram_renable;
  wire [32-1:0] _mul_5_y_source_ram_rdata;
  reg _mul_5_y_source_fifo_deq;
  wire [32-1:0] _mul_5_y_source_fifo_rdata;
  reg [32-1:0] _mul_5_y_source_empty_data;
  reg _mul_5_rshift_idle;
  reg [33-1:0] _mul_5_rshift_source_count;
  reg [5-1:0] _mul_5_rshift_source_mode;
  reg [16-1:0] _mul_5_rshift_source_generator_id;
  reg [32-1:0] _mul_5_rshift_source_offset;
  reg [33-1:0] _mul_5_rshift_source_size;
  reg [32-1:0] _mul_5_rshift_source_stride;
  reg [32-1:0] _mul_5_rshift_source_offset_buf;
  reg [33-1:0] _mul_5_rshift_source_size_buf;
  reg [32-1:0] _mul_5_rshift_source_stride_buf;
  reg [8-1:0] _mul_5_rshift_source_sel;
  reg [32-1:0] _mul_5_rshift_source_ram_raddr;
  reg _mul_5_rshift_source_ram_renable;
  wire [32-1:0] _mul_5_rshift_source_ram_rdata;
  reg _mul_5_rshift_source_fifo_deq;
  wire [32-1:0] _mul_5_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_5_rshift_source_empty_data;
  reg [33-1:0] _mul_5_z_sink_count;
  reg [5-1:0] _mul_5_z_sink_mode;
  reg [16-1:0] _mul_5_z_sink_generator_id;
  reg [32-1:0] _mul_5_z_sink_offset;
  reg [33-1:0] _mul_5_z_sink_size;
  reg [32-1:0] _mul_5_z_sink_stride;
  reg [32-1:0] _mul_5_z_sink_offset_buf;
  reg [33-1:0] _mul_5_z_sink_size_buf;
  reg [32-1:0] _mul_5_z_sink_stride_buf;
  reg [8-1:0] _mul_5_z_sink_sel;
  reg [32-1:0] _mul_5_z_sink_waddr;
  reg _mul_5_z_sink_wenable;
  reg [64-1:0] _mul_5_z_sink_wdata;
  reg _mul_5_z_sink_fifo_enq;
  reg [64-1:0] _mul_5_z_sink_fifo_wdata;
  reg [64-1:0] _mul_5_z_sink_immediate;
  reg _mul_6_stream_ivalid;
  wire _mul_6_stream_oready;
  wire _mul_6_stream_internal_oready;
  assign _mul_6_stream_internal_oready = 1;
  reg [32-1:0] _mul_6_fsm;
  localparam _mul_6_fsm_init = 0;
  wire _mul_6_run_flag;
  assign _mul_6_run_flag = 0;
  reg _mul_6_source_start;
  wire _mul_6_source_stop;
  reg _mul_6_source_busy;
  wire _mul_6_sink_start;
  wire _mul_6_sink_stop;
  wire _mul_6_sink_busy;
  wire _mul_6_busy;
  reg _mul_6_busy_reg;
  wire _mul_6_is_root;
  reg _mul_6_x_idle;
  reg [33-1:0] _mul_6_x_source_count;
  reg [5-1:0] _mul_6_x_source_mode;
  reg [16-1:0] _mul_6_x_source_generator_id;
  reg [32-1:0] _mul_6_x_source_offset;
  reg [33-1:0] _mul_6_x_source_size;
  reg [32-1:0] _mul_6_x_source_stride;
  reg [32-1:0] _mul_6_x_source_offset_buf;
  reg [33-1:0] _mul_6_x_source_size_buf;
  reg [32-1:0] _mul_6_x_source_stride_buf;
  reg [8-1:0] _mul_6_x_source_sel;
  reg [32-1:0] _mul_6_x_source_ram_raddr;
  reg _mul_6_x_source_ram_renable;
  wire [32-1:0] _mul_6_x_source_ram_rdata;
  reg _mul_6_x_source_fifo_deq;
  wire [32-1:0] _mul_6_x_source_fifo_rdata;
  reg [32-1:0] _mul_6_x_source_empty_data;
  reg _mul_6_y_idle;
  reg [33-1:0] _mul_6_y_source_count;
  reg [5-1:0] _mul_6_y_source_mode;
  reg [16-1:0] _mul_6_y_source_generator_id;
  reg [32-1:0] _mul_6_y_source_offset;
  reg [33-1:0] _mul_6_y_source_size;
  reg [32-1:0] _mul_6_y_source_stride;
  reg [32-1:0] _mul_6_y_source_offset_buf;
  reg [33-1:0] _mul_6_y_source_size_buf;
  reg [32-1:0] _mul_6_y_source_stride_buf;
  reg [8-1:0] _mul_6_y_source_sel;
  reg [32-1:0] _mul_6_y_source_ram_raddr;
  reg _mul_6_y_source_ram_renable;
  wire [32-1:0] _mul_6_y_source_ram_rdata;
  reg _mul_6_y_source_fifo_deq;
  wire [32-1:0] _mul_6_y_source_fifo_rdata;
  reg [32-1:0] _mul_6_y_source_empty_data;
  reg _mul_6_rshift_idle;
  reg [33-1:0] _mul_6_rshift_source_count;
  reg [5-1:0] _mul_6_rshift_source_mode;
  reg [16-1:0] _mul_6_rshift_source_generator_id;
  reg [32-1:0] _mul_6_rshift_source_offset;
  reg [33-1:0] _mul_6_rshift_source_size;
  reg [32-1:0] _mul_6_rshift_source_stride;
  reg [32-1:0] _mul_6_rshift_source_offset_buf;
  reg [33-1:0] _mul_6_rshift_source_size_buf;
  reg [32-1:0] _mul_6_rshift_source_stride_buf;
  reg [8-1:0] _mul_6_rshift_source_sel;
  reg [32-1:0] _mul_6_rshift_source_ram_raddr;
  reg _mul_6_rshift_source_ram_renable;
  wire [32-1:0] _mul_6_rshift_source_ram_rdata;
  reg _mul_6_rshift_source_fifo_deq;
  wire [32-1:0] _mul_6_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_6_rshift_source_empty_data;
  reg [33-1:0] _mul_6_z_sink_count;
  reg [5-1:0] _mul_6_z_sink_mode;
  reg [16-1:0] _mul_6_z_sink_generator_id;
  reg [32-1:0] _mul_6_z_sink_offset;
  reg [33-1:0] _mul_6_z_sink_size;
  reg [32-1:0] _mul_6_z_sink_stride;
  reg [32-1:0] _mul_6_z_sink_offset_buf;
  reg [33-1:0] _mul_6_z_sink_size_buf;
  reg [32-1:0] _mul_6_z_sink_stride_buf;
  reg [8-1:0] _mul_6_z_sink_sel;
  reg [32-1:0] _mul_6_z_sink_waddr;
  reg _mul_6_z_sink_wenable;
  reg [64-1:0] _mul_6_z_sink_wdata;
  reg _mul_6_z_sink_fifo_enq;
  reg [64-1:0] _mul_6_z_sink_fifo_wdata;
  reg [64-1:0] _mul_6_z_sink_immediate;
  reg _mul_7_stream_ivalid;
  wire _mul_7_stream_oready;
  wire _mul_7_stream_internal_oready;
  assign _mul_7_stream_internal_oready = 1;
  reg [32-1:0] _mul_7_fsm;
  localparam _mul_7_fsm_init = 0;
  wire _mul_7_run_flag;
  assign _mul_7_run_flag = 0;
  reg _mul_7_source_start;
  wire _mul_7_source_stop;
  reg _mul_7_source_busy;
  wire _mul_7_sink_start;
  wire _mul_7_sink_stop;
  wire _mul_7_sink_busy;
  wire _mul_7_busy;
  reg _mul_7_busy_reg;
  wire _mul_7_is_root;
  reg _mul_7_x_idle;
  reg [33-1:0] _mul_7_x_source_count;
  reg [5-1:0] _mul_7_x_source_mode;
  reg [16-1:0] _mul_7_x_source_generator_id;
  reg [32-1:0] _mul_7_x_source_offset;
  reg [33-1:0] _mul_7_x_source_size;
  reg [32-1:0] _mul_7_x_source_stride;
  reg [32-1:0] _mul_7_x_source_offset_buf;
  reg [33-1:0] _mul_7_x_source_size_buf;
  reg [32-1:0] _mul_7_x_source_stride_buf;
  reg [8-1:0] _mul_7_x_source_sel;
  reg [32-1:0] _mul_7_x_source_ram_raddr;
  reg _mul_7_x_source_ram_renable;
  wire [32-1:0] _mul_7_x_source_ram_rdata;
  reg _mul_7_x_source_fifo_deq;
  wire [32-1:0] _mul_7_x_source_fifo_rdata;
  reg [32-1:0] _mul_7_x_source_empty_data;
  reg _mul_7_y_idle;
  reg [33-1:0] _mul_7_y_source_count;
  reg [5-1:0] _mul_7_y_source_mode;
  reg [16-1:0] _mul_7_y_source_generator_id;
  reg [32-1:0] _mul_7_y_source_offset;
  reg [33-1:0] _mul_7_y_source_size;
  reg [32-1:0] _mul_7_y_source_stride;
  reg [32-1:0] _mul_7_y_source_offset_buf;
  reg [33-1:0] _mul_7_y_source_size_buf;
  reg [32-1:0] _mul_7_y_source_stride_buf;
  reg [8-1:0] _mul_7_y_source_sel;
  reg [32-1:0] _mul_7_y_source_ram_raddr;
  reg _mul_7_y_source_ram_renable;
  wire [32-1:0] _mul_7_y_source_ram_rdata;
  reg _mul_7_y_source_fifo_deq;
  wire [32-1:0] _mul_7_y_source_fifo_rdata;
  reg [32-1:0] _mul_7_y_source_empty_data;
  reg _mul_7_rshift_idle;
  reg [33-1:0] _mul_7_rshift_source_count;
  reg [5-1:0] _mul_7_rshift_source_mode;
  reg [16-1:0] _mul_7_rshift_source_generator_id;
  reg [32-1:0] _mul_7_rshift_source_offset;
  reg [33-1:0] _mul_7_rshift_source_size;
  reg [32-1:0] _mul_7_rshift_source_stride;
  reg [32-1:0] _mul_7_rshift_source_offset_buf;
  reg [33-1:0] _mul_7_rshift_source_size_buf;
  reg [32-1:0] _mul_7_rshift_source_stride_buf;
  reg [8-1:0] _mul_7_rshift_source_sel;
  reg [32-1:0] _mul_7_rshift_source_ram_raddr;
  reg _mul_7_rshift_source_ram_renable;
  wire [32-1:0] _mul_7_rshift_source_ram_rdata;
  reg _mul_7_rshift_source_fifo_deq;
  wire [32-1:0] _mul_7_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_7_rshift_source_empty_data;
  reg [33-1:0] _mul_7_z_sink_count;
  reg [5-1:0] _mul_7_z_sink_mode;
  reg [16-1:0] _mul_7_z_sink_generator_id;
  reg [32-1:0] _mul_7_z_sink_offset;
  reg [33-1:0] _mul_7_z_sink_size;
  reg [32-1:0] _mul_7_z_sink_stride;
  reg [32-1:0] _mul_7_z_sink_offset_buf;
  reg [33-1:0] _mul_7_z_sink_size_buf;
  reg [32-1:0] _mul_7_z_sink_stride_buf;
  reg [8-1:0] _mul_7_z_sink_sel;
  reg [32-1:0] _mul_7_z_sink_waddr;
  reg _mul_7_z_sink_wenable;
  reg [64-1:0] _mul_7_z_sink_wdata;
  reg _mul_7_z_sink_fifo_enq;
  reg [64-1:0] _mul_7_z_sink_fifo_wdata;
  reg [64-1:0] _mul_7_z_sink_immediate;
  reg _mul_8_stream_ivalid;
  wire _mul_8_stream_oready;
  wire _mul_8_stream_internal_oready;
  assign _mul_8_stream_internal_oready = 1;
  reg [32-1:0] _mul_8_fsm;
  localparam _mul_8_fsm_init = 0;
  wire _mul_8_run_flag;
  assign _mul_8_run_flag = 0;
  reg _mul_8_source_start;
  wire _mul_8_source_stop;
  reg _mul_8_source_busy;
  wire _mul_8_sink_start;
  wire _mul_8_sink_stop;
  wire _mul_8_sink_busy;
  wire _mul_8_busy;
  reg _mul_8_busy_reg;
  wire _mul_8_is_root;
  reg _mul_8_x_idle;
  reg [33-1:0] _mul_8_x_source_count;
  reg [5-1:0] _mul_8_x_source_mode;
  reg [16-1:0] _mul_8_x_source_generator_id;
  reg [32-1:0] _mul_8_x_source_offset;
  reg [33-1:0] _mul_8_x_source_size;
  reg [32-1:0] _mul_8_x_source_stride;
  reg [32-1:0] _mul_8_x_source_offset_buf;
  reg [33-1:0] _mul_8_x_source_size_buf;
  reg [32-1:0] _mul_8_x_source_stride_buf;
  reg [8-1:0] _mul_8_x_source_sel;
  reg [32-1:0] _mul_8_x_source_ram_raddr;
  reg _mul_8_x_source_ram_renable;
  wire [32-1:0] _mul_8_x_source_ram_rdata;
  reg _mul_8_x_source_fifo_deq;
  wire [32-1:0] _mul_8_x_source_fifo_rdata;
  reg [32-1:0] _mul_8_x_source_empty_data;
  reg _mul_8_y_idle;
  reg [33-1:0] _mul_8_y_source_count;
  reg [5-1:0] _mul_8_y_source_mode;
  reg [16-1:0] _mul_8_y_source_generator_id;
  reg [32-1:0] _mul_8_y_source_offset;
  reg [33-1:0] _mul_8_y_source_size;
  reg [32-1:0] _mul_8_y_source_stride;
  reg [32-1:0] _mul_8_y_source_offset_buf;
  reg [33-1:0] _mul_8_y_source_size_buf;
  reg [32-1:0] _mul_8_y_source_stride_buf;
  reg [8-1:0] _mul_8_y_source_sel;
  reg [32-1:0] _mul_8_y_source_ram_raddr;
  reg _mul_8_y_source_ram_renable;
  wire [32-1:0] _mul_8_y_source_ram_rdata;
  reg _mul_8_y_source_fifo_deq;
  wire [32-1:0] _mul_8_y_source_fifo_rdata;
  reg [32-1:0] _mul_8_y_source_empty_data;
  reg _mul_8_rshift_idle;
  reg [33-1:0] _mul_8_rshift_source_count;
  reg [5-1:0] _mul_8_rshift_source_mode;
  reg [16-1:0] _mul_8_rshift_source_generator_id;
  reg [32-1:0] _mul_8_rshift_source_offset;
  reg [33-1:0] _mul_8_rshift_source_size;
  reg [32-1:0] _mul_8_rshift_source_stride;
  reg [32-1:0] _mul_8_rshift_source_offset_buf;
  reg [33-1:0] _mul_8_rshift_source_size_buf;
  reg [32-1:0] _mul_8_rshift_source_stride_buf;
  reg [8-1:0] _mul_8_rshift_source_sel;
  reg [32-1:0] _mul_8_rshift_source_ram_raddr;
  reg _mul_8_rshift_source_ram_renable;
  wire [32-1:0] _mul_8_rshift_source_ram_rdata;
  reg _mul_8_rshift_source_fifo_deq;
  wire [32-1:0] _mul_8_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_8_rshift_source_empty_data;
  reg [33-1:0] _mul_8_z_sink_count;
  reg [5-1:0] _mul_8_z_sink_mode;
  reg [16-1:0] _mul_8_z_sink_generator_id;
  reg [32-1:0] _mul_8_z_sink_offset;
  reg [33-1:0] _mul_8_z_sink_size;
  reg [32-1:0] _mul_8_z_sink_stride;
  reg [32-1:0] _mul_8_z_sink_offset_buf;
  reg [33-1:0] _mul_8_z_sink_size_buf;
  reg [32-1:0] _mul_8_z_sink_stride_buf;
  reg [8-1:0] _mul_8_z_sink_sel;
  reg [32-1:0] _mul_8_z_sink_waddr;
  reg _mul_8_z_sink_wenable;
  reg [64-1:0] _mul_8_z_sink_wdata;
  reg _mul_8_z_sink_fifo_enq;
  reg [64-1:0] _mul_8_z_sink_fifo_wdata;
  reg [64-1:0] _mul_8_z_sink_immediate;
  reg _mul_9_stream_ivalid;
  wire _mul_9_stream_oready;
  wire _mul_9_stream_internal_oready;
  assign _mul_9_stream_internal_oready = 1;
  reg [32-1:0] _mul_9_fsm;
  localparam _mul_9_fsm_init = 0;
  wire _mul_9_run_flag;
  assign _mul_9_run_flag = 0;
  reg _mul_9_source_start;
  wire _mul_9_source_stop;
  reg _mul_9_source_busy;
  wire _mul_9_sink_start;
  wire _mul_9_sink_stop;
  wire _mul_9_sink_busy;
  wire _mul_9_busy;
  reg _mul_9_busy_reg;
  wire _mul_9_is_root;
  reg _mul_9_x_idle;
  reg [33-1:0] _mul_9_x_source_count;
  reg [5-1:0] _mul_9_x_source_mode;
  reg [16-1:0] _mul_9_x_source_generator_id;
  reg [32-1:0] _mul_9_x_source_offset;
  reg [33-1:0] _mul_9_x_source_size;
  reg [32-1:0] _mul_9_x_source_stride;
  reg [32-1:0] _mul_9_x_source_offset_buf;
  reg [33-1:0] _mul_9_x_source_size_buf;
  reg [32-1:0] _mul_9_x_source_stride_buf;
  reg [8-1:0] _mul_9_x_source_sel;
  reg [32-1:0] _mul_9_x_source_ram_raddr;
  reg _mul_9_x_source_ram_renable;
  wire [32-1:0] _mul_9_x_source_ram_rdata;
  reg _mul_9_x_source_fifo_deq;
  wire [32-1:0] _mul_9_x_source_fifo_rdata;
  reg [32-1:0] _mul_9_x_source_empty_data;
  reg _mul_9_y_idle;
  reg [33-1:0] _mul_9_y_source_count;
  reg [5-1:0] _mul_9_y_source_mode;
  reg [16-1:0] _mul_9_y_source_generator_id;
  reg [32-1:0] _mul_9_y_source_offset;
  reg [33-1:0] _mul_9_y_source_size;
  reg [32-1:0] _mul_9_y_source_stride;
  reg [32-1:0] _mul_9_y_source_offset_buf;
  reg [33-1:0] _mul_9_y_source_size_buf;
  reg [32-1:0] _mul_9_y_source_stride_buf;
  reg [8-1:0] _mul_9_y_source_sel;
  reg [32-1:0] _mul_9_y_source_ram_raddr;
  reg _mul_9_y_source_ram_renable;
  wire [32-1:0] _mul_9_y_source_ram_rdata;
  reg _mul_9_y_source_fifo_deq;
  wire [32-1:0] _mul_9_y_source_fifo_rdata;
  reg [32-1:0] _mul_9_y_source_empty_data;
  reg _mul_9_rshift_idle;
  reg [33-1:0] _mul_9_rshift_source_count;
  reg [5-1:0] _mul_9_rshift_source_mode;
  reg [16-1:0] _mul_9_rshift_source_generator_id;
  reg [32-1:0] _mul_9_rshift_source_offset;
  reg [33-1:0] _mul_9_rshift_source_size;
  reg [32-1:0] _mul_9_rshift_source_stride;
  reg [32-1:0] _mul_9_rshift_source_offset_buf;
  reg [33-1:0] _mul_9_rshift_source_size_buf;
  reg [32-1:0] _mul_9_rshift_source_stride_buf;
  reg [8-1:0] _mul_9_rshift_source_sel;
  reg [32-1:0] _mul_9_rshift_source_ram_raddr;
  reg _mul_9_rshift_source_ram_renable;
  wire [32-1:0] _mul_9_rshift_source_ram_rdata;
  reg _mul_9_rshift_source_fifo_deq;
  wire [32-1:0] _mul_9_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_9_rshift_source_empty_data;
  reg [33-1:0] _mul_9_z_sink_count;
  reg [5-1:0] _mul_9_z_sink_mode;
  reg [16-1:0] _mul_9_z_sink_generator_id;
  reg [32-1:0] _mul_9_z_sink_offset;
  reg [33-1:0] _mul_9_z_sink_size;
  reg [32-1:0] _mul_9_z_sink_stride;
  reg [32-1:0] _mul_9_z_sink_offset_buf;
  reg [33-1:0] _mul_9_z_sink_size_buf;
  reg [32-1:0] _mul_9_z_sink_stride_buf;
  reg [8-1:0] _mul_9_z_sink_sel;
  reg [32-1:0] _mul_9_z_sink_waddr;
  reg _mul_9_z_sink_wenable;
  reg [64-1:0] _mul_9_z_sink_wdata;
  reg _mul_9_z_sink_fifo_enq;
  reg [64-1:0] _mul_9_z_sink_fifo_wdata;
  reg [64-1:0] _mul_9_z_sink_immediate;
  reg _mul_10_stream_ivalid;
  wire _mul_10_stream_oready;
  wire _mul_10_stream_internal_oready;
  assign _mul_10_stream_internal_oready = 1;
  reg [32-1:0] _mul_10_fsm;
  localparam _mul_10_fsm_init = 0;
  wire _mul_10_run_flag;
  assign _mul_10_run_flag = 0;
  reg _mul_10_source_start;
  wire _mul_10_source_stop;
  reg _mul_10_source_busy;
  wire _mul_10_sink_start;
  wire _mul_10_sink_stop;
  wire _mul_10_sink_busy;
  wire _mul_10_busy;
  reg _mul_10_busy_reg;
  wire _mul_10_is_root;
  reg _mul_10_x_idle;
  reg [33-1:0] _mul_10_x_source_count;
  reg [5-1:0] _mul_10_x_source_mode;
  reg [16-1:0] _mul_10_x_source_generator_id;
  reg [32-1:0] _mul_10_x_source_offset;
  reg [33-1:0] _mul_10_x_source_size;
  reg [32-1:0] _mul_10_x_source_stride;
  reg [32-1:0] _mul_10_x_source_offset_buf;
  reg [33-1:0] _mul_10_x_source_size_buf;
  reg [32-1:0] _mul_10_x_source_stride_buf;
  reg [8-1:0] _mul_10_x_source_sel;
  reg [32-1:0] _mul_10_x_source_ram_raddr;
  reg _mul_10_x_source_ram_renable;
  wire [32-1:0] _mul_10_x_source_ram_rdata;
  reg _mul_10_x_source_fifo_deq;
  wire [32-1:0] _mul_10_x_source_fifo_rdata;
  reg [32-1:0] _mul_10_x_source_empty_data;
  reg _mul_10_y_idle;
  reg [33-1:0] _mul_10_y_source_count;
  reg [5-1:0] _mul_10_y_source_mode;
  reg [16-1:0] _mul_10_y_source_generator_id;
  reg [32-1:0] _mul_10_y_source_offset;
  reg [33-1:0] _mul_10_y_source_size;
  reg [32-1:0] _mul_10_y_source_stride;
  reg [32-1:0] _mul_10_y_source_offset_buf;
  reg [33-1:0] _mul_10_y_source_size_buf;
  reg [32-1:0] _mul_10_y_source_stride_buf;
  reg [8-1:0] _mul_10_y_source_sel;
  reg [32-1:0] _mul_10_y_source_ram_raddr;
  reg _mul_10_y_source_ram_renable;
  wire [32-1:0] _mul_10_y_source_ram_rdata;
  reg _mul_10_y_source_fifo_deq;
  wire [32-1:0] _mul_10_y_source_fifo_rdata;
  reg [32-1:0] _mul_10_y_source_empty_data;
  reg _mul_10_rshift_idle;
  reg [33-1:0] _mul_10_rshift_source_count;
  reg [5-1:0] _mul_10_rshift_source_mode;
  reg [16-1:0] _mul_10_rshift_source_generator_id;
  reg [32-1:0] _mul_10_rshift_source_offset;
  reg [33-1:0] _mul_10_rshift_source_size;
  reg [32-1:0] _mul_10_rshift_source_stride;
  reg [32-1:0] _mul_10_rshift_source_offset_buf;
  reg [33-1:0] _mul_10_rshift_source_size_buf;
  reg [32-1:0] _mul_10_rshift_source_stride_buf;
  reg [8-1:0] _mul_10_rshift_source_sel;
  reg [32-1:0] _mul_10_rshift_source_ram_raddr;
  reg _mul_10_rshift_source_ram_renable;
  wire [32-1:0] _mul_10_rshift_source_ram_rdata;
  reg _mul_10_rshift_source_fifo_deq;
  wire [32-1:0] _mul_10_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_10_rshift_source_empty_data;
  reg [33-1:0] _mul_10_z_sink_count;
  reg [5-1:0] _mul_10_z_sink_mode;
  reg [16-1:0] _mul_10_z_sink_generator_id;
  reg [32-1:0] _mul_10_z_sink_offset;
  reg [33-1:0] _mul_10_z_sink_size;
  reg [32-1:0] _mul_10_z_sink_stride;
  reg [32-1:0] _mul_10_z_sink_offset_buf;
  reg [33-1:0] _mul_10_z_sink_size_buf;
  reg [32-1:0] _mul_10_z_sink_stride_buf;
  reg [8-1:0] _mul_10_z_sink_sel;
  reg [32-1:0] _mul_10_z_sink_waddr;
  reg _mul_10_z_sink_wenable;
  reg [64-1:0] _mul_10_z_sink_wdata;
  reg _mul_10_z_sink_fifo_enq;
  reg [64-1:0] _mul_10_z_sink_fifo_wdata;
  reg [64-1:0] _mul_10_z_sink_immediate;
  reg _mul_11_stream_ivalid;
  wire _mul_11_stream_oready;
  wire _mul_11_stream_internal_oready;
  assign _mul_11_stream_internal_oready = 1;
  reg [32-1:0] _mul_11_fsm;
  localparam _mul_11_fsm_init = 0;
  wire _mul_11_run_flag;
  assign _mul_11_run_flag = 0;
  reg _mul_11_source_start;
  wire _mul_11_source_stop;
  reg _mul_11_source_busy;
  wire _mul_11_sink_start;
  wire _mul_11_sink_stop;
  wire _mul_11_sink_busy;
  wire _mul_11_busy;
  reg _mul_11_busy_reg;
  wire _mul_11_is_root;
  reg _mul_11_x_idle;
  reg [33-1:0] _mul_11_x_source_count;
  reg [5-1:0] _mul_11_x_source_mode;
  reg [16-1:0] _mul_11_x_source_generator_id;
  reg [32-1:0] _mul_11_x_source_offset;
  reg [33-1:0] _mul_11_x_source_size;
  reg [32-1:0] _mul_11_x_source_stride;
  reg [32-1:0] _mul_11_x_source_offset_buf;
  reg [33-1:0] _mul_11_x_source_size_buf;
  reg [32-1:0] _mul_11_x_source_stride_buf;
  reg [8-1:0] _mul_11_x_source_sel;
  reg [32-1:0] _mul_11_x_source_ram_raddr;
  reg _mul_11_x_source_ram_renable;
  wire [32-1:0] _mul_11_x_source_ram_rdata;
  reg _mul_11_x_source_fifo_deq;
  wire [32-1:0] _mul_11_x_source_fifo_rdata;
  reg [32-1:0] _mul_11_x_source_empty_data;
  reg _mul_11_y_idle;
  reg [33-1:0] _mul_11_y_source_count;
  reg [5-1:0] _mul_11_y_source_mode;
  reg [16-1:0] _mul_11_y_source_generator_id;
  reg [32-1:0] _mul_11_y_source_offset;
  reg [33-1:0] _mul_11_y_source_size;
  reg [32-1:0] _mul_11_y_source_stride;
  reg [32-1:0] _mul_11_y_source_offset_buf;
  reg [33-1:0] _mul_11_y_source_size_buf;
  reg [32-1:0] _mul_11_y_source_stride_buf;
  reg [8-1:0] _mul_11_y_source_sel;
  reg [32-1:0] _mul_11_y_source_ram_raddr;
  reg _mul_11_y_source_ram_renable;
  wire [32-1:0] _mul_11_y_source_ram_rdata;
  reg _mul_11_y_source_fifo_deq;
  wire [32-1:0] _mul_11_y_source_fifo_rdata;
  reg [32-1:0] _mul_11_y_source_empty_data;
  reg _mul_11_rshift_idle;
  reg [33-1:0] _mul_11_rshift_source_count;
  reg [5-1:0] _mul_11_rshift_source_mode;
  reg [16-1:0] _mul_11_rshift_source_generator_id;
  reg [32-1:0] _mul_11_rshift_source_offset;
  reg [33-1:0] _mul_11_rshift_source_size;
  reg [32-1:0] _mul_11_rshift_source_stride;
  reg [32-1:0] _mul_11_rshift_source_offset_buf;
  reg [33-1:0] _mul_11_rshift_source_size_buf;
  reg [32-1:0] _mul_11_rshift_source_stride_buf;
  reg [8-1:0] _mul_11_rshift_source_sel;
  reg [32-1:0] _mul_11_rshift_source_ram_raddr;
  reg _mul_11_rshift_source_ram_renable;
  wire [32-1:0] _mul_11_rshift_source_ram_rdata;
  reg _mul_11_rshift_source_fifo_deq;
  wire [32-1:0] _mul_11_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_11_rshift_source_empty_data;
  reg [33-1:0] _mul_11_z_sink_count;
  reg [5-1:0] _mul_11_z_sink_mode;
  reg [16-1:0] _mul_11_z_sink_generator_id;
  reg [32-1:0] _mul_11_z_sink_offset;
  reg [33-1:0] _mul_11_z_sink_size;
  reg [32-1:0] _mul_11_z_sink_stride;
  reg [32-1:0] _mul_11_z_sink_offset_buf;
  reg [33-1:0] _mul_11_z_sink_size_buf;
  reg [32-1:0] _mul_11_z_sink_stride_buf;
  reg [8-1:0] _mul_11_z_sink_sel;
  reg [32-1:0] _mul_11_z_sink_waddr;
  reg _mul_11_z_sink_wenable;
  reg [64-1:0] _mul_11_z_sink_wdata;
  reg _mul_11_z_sink_fifo_enq;
  reg [64-1:0] _mul_11_z_sink_fifo_wdata;
  reg [64-1:0] _mul_11_z_sink_immediate;
  reg _mul_12_stream_ivalid;
  wire _mul_12_stream_oready;
  wire _mul_12_stream_internal_oready;
  assign _mul_12_stream_internal_oready = 1;
  reg [32-1:0] _mul_12_fsm;
  localparam _mul_12_fsm_init = 0;
  wire _mul_12_run_flag;
  assign _mul_12_run_flag = 0;
  reg _mul_12_source_start;
  wire _mul_12_source_stop;
  reg _mul_12_source_busy;
  wire _mul_12_sink_start;
  wire _mul_12_sink_stop;
  wire _mul_12_sink_busy;
  wire _mul_12_busy;
  reg _mul_12_busy_reg;
  wire _mul_12_is_root;
  reg _mul_12_x_idle;
  reg [33-1:0] _mul_12_x_source_count;
  reg [5-1:0] _mul_12_x_source_mode;
  reg [16-1:0] _mul_12_x_source_generator_id;
  reg [32-1:0] _mul_12_x_source_offset;
  reg [33-1:0] _mul_12_x_source_size;
  reg [32-1:0] _mul_12_x_source_stride;
  reg [32-1:0] _mul_12_x_source_offset_buf;
  reg [33-1:0] _mul_12_x_source_size_buf;
  reg [32-1:0] _mul_12_x_source_stride_buf;
  reg [8-1:0] _mul_12_x_source_sel;
  reg [32-1:0] _mul_12_x_source_ram_raddr;
  reg _mul_12_x_source_ram_renable;
  wire [32-1:0] _mul_12_x_source_ram_rdata;
  reg _mul_12_x_source_fifo_deq;
  wire [32-1:0] _mul_12_x_source_fifo_rdata;
  reg [32-1:0] _mul_12_x_source_empty_data;
  reg _mul_12_y_idle;
  reg [33-1:0] _mul_12_y_source_count;
  reg [5-1:0] _mul_12_y_source_mode;
  reg [16-1:0] _mul_12_y_source_generator_id;
  reg [32-1:0] _mul_12_y_source_offset;
  reg [33-1:0] _mul_12_y_source_size;
  reg [32-1:0] _mul_12_y_source_stride;
  reg [32-1:0] _mul_12_y_source_offset_buf;
  reg [33-1:0] _mul_12_y_source_size_buf;
  reg [32-1:0] _mul_12_y_source_stride_buf;
  reg [8-1:0] _mul_12_y_source_sel;
  reg [32-1:0] _mul_12_y_source_ram_raddr;
  reg _mul_12_y_source_ram_renable;
  wire [32-1:0] _mul_12_y_source_ram_rdata;
  reg _mul_12_y_source_fifo_deq;
  wire [32-1:0] _mul_12_y_source_fifo_rdata;
  reg [32-1:0] _mul_12_y_source_empty_data;
  reg _mul_12_rshift_idle;
  reg [33-1:0] _mul_12_rshift_source_count;
  reg [5-1:0] _mul_12_rshift_source_mode;
  reg [16-1:0] _mul_12_rshift_source_generator_id;
  reg [32-1:0] _mul_12_rshift_source_offset;
  reg [33-1:0] _mul_12_rshift_source_size;
  reg [32-1:0] _mul_12_rshift_source_stride;
  reg [32-1:0] _mul_12_rshift_source_offset_buf;
  reg [33-1:0] _mul_12_rshift_source_size_buf;
  reg [32-1:0] _mul_12_rshift_source_stride_buf;
  reg [8-1:0] _mul_12_rshift_source_sel;
  reg [32-1:0] _mul_12_rshift_source_ram_raddr;
  reg _mul_12_rshift_source_ram_renable;
  wire [32-1:0] _mul_12_rshift_source_ram_rdata;
  reg _mul_12_rshift_source_fifo_deq;
  wire [32-1:0] _mul_12_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_12_rshift_source_empty_data;
  reg [33-1:0] _mul_12_z_sink_count;
  reg [5-1:0] _mul_12_z_sink_mode;
  reg [16-1:0] _mul_12_z_sink_generator_id;
  reg [32-1:0] _mul_12_z_sink_offset;
  reg [33-1:0] _mul_12_z_sink_size;
  reg [32-1:0] _mul_12_z_sink_stride;
  reg [32-1:0] _mul_12_z_sink_offset_buf;
  reg [33-1:0] _mul_12_z_sink_size_buf;
  reg [32-1:0] _mul_12_z_sink_stride_buf;
  reg [8-1:0] _mul_12_z_sink_sel;
  reg [32-1:0] _mul_12_z_sink_waddr;
  reg _mul_12_z_sink_wenable;
  reg [64-1:0] _mul_12_z_sink_wdata;
  reg _mul_12_z_sink_fifo_enq;
  reg [64-1:0] _mul_12_z_sink_fifo_wdata;
  reg [64-1:0] _mul_12_z_sink_immediate;
  reg __reduce_max_13_stream_ivalid;
  wire __reduce_max_13_stream_oready;
  wire __reduce_max_13_stream_internal_oready;
  assign __reduce_max_13_stream_internal_oready = 1;
  reg [32-1:0] __reduce_max_13_fsm;
  localparam __reduce_max_13_fsm_init = 0;
  wire __reduce_max_13_run_flag;
  assign __reduce_max_13_run_flag = 0;
  reg __reduce_max_13_source_start;
  wire __reduce_max_13_source_stop;
  reg __reduce_max_13_source_busy;
  wire __reduce_max_13_sink_start;
  wire __reduce_max_13_sink_stop;
  wire __reduce_max_13_sink_busy;
  wire __reduce_max_13_busy;
  reg __reduce_max_13_busy_reg;
  wire __reduce_max_13_is_root;
  reg __reduce_max_13_x_idle;
  reg [33-1:0] __reduce_max_13_x_source_count;
  reg [5-1:0] __reduce_max_13_x_source_mode;
  reg [16-1:0] __reduce_max_13_x_source_generator_id;
  reg [32-1:0] __reduce_max_13_x_source_offset;
  reg [33-1:0] __reduce_max_13_x_source_size;
  reg [32-1:0] __reduce_max_13_x_source_stride;
  reg [32-1:0] __reduce_max_13_x_source_offset_buf;
  reg [33-1:0] __reduce_max_13_x_source_size_buf;
  reg [32-1:0] __reduce_max_13_x_source_stride_buf;
  reg [8-1:0] __reduce_max_13_x_source_sel;
  reg [32-1:0] __reduce_max_13_x_source_ram_raddr;
  reg __reduce_max_13_x_source_ram_renable;
  wire [32-1:0] __reduce_max_13_x_source_ram_rdata;
  reg __reduce_max_13_x_source_fifo_deq;
  wire [32-1:0] __reduce_max_13_x_source_fifo_rdata;
  reg [32-1:0] __reduce_max_13_x_source_empty_data;
  reg [32-1:0] __reduce_max_13_size_next_parameter_data;
  reg [33-1:0] __reduce_max_13_data_sink_count;
  reg [5-1:0] __reduce_max_13_data_sink_mode;
  reg [16-1:0] __reduce_max_13_data_sink_generator_id;
  reg [32-1:0] __reduce_max_13_data_sink_offset;
  reg [33-1:0] __reduce_max_13_data_sink_size;
  reg [32-1:0] __reduce_max_13_data_sink_stride;
  reg [32-1:0] __reduce_max_13_data_sink_offset_buf;
  reg [33-1:0] __reduce_max_13_data_sink_size_buf;
  reg [32-1:0] __reduce_max_13_data_sink_stride_buf;
  reg [8-1:0] __reduce_max_13_data_sink_sel;
  reg [32-1:0] __reduce_max_13_data_sink_waddr;
  reg __reduce_max_13_data_sink_wenable;
  reg [32-1:0] __reduce_max_13_data_sink_wdata;
  reg __reduce_max_13_data_sink_fifo_enq;
  reg [32-1:0] __reduce_max_13_data_sink_fifo_wdata;
  reg [32-1:0] __reduce_max_13_data_sink_immediate;
  reg [33-1:0] __reduce_max_13_valid_sink_count;
  reg [5-1:0] __reduce_max_13_valid_sink_mode;
  reg [16-1:0] __reduce_max_13_valid_sink_generator_id;
  reg [32-1:0] __reduce_max_13_valid_sink_offset;
  reg [33-1:0] __reduce_max_13_valid_sink_size;
  reg [32-1:0] __reduce_max_13_valid_sink_stride;
  reg [32-1:0] __reduce_max_13_valid_sink_offset_buf;
  reg [33-1:0] __reduce_max_13_valid_sink_size_buf;
  reg [32-1:0] __reduce_max_13_valid_sink_stride_buf;
  reg [8-1:0] __reduce_max_13_valid_sink_sel;
  reg [32-1:0] __reduce_max_13_valid_sink_waddr;
  reg __reduce_max_13_valid_sink_wenable;
  reg [1-1:0] __reduce_max_13_valid_sink_wdata;
  reg __reduce_max_13_valid_sink_fifo_enq;
  reg [1-1:0] __reduce_max_13_valid_sink_fifo_wdata;
  reg [1-1:0] __reduce_max_13_valid_sink_immediate;
  reg _stream_conv2d_25_stream_ivalid;
  wire _stream_conv2d_25_stream_oready;
  wire _stream_conv2d_25_stream_internal_oready;
  assign _stream_conv2d_25_stream_oready = _stream_conv2d_25_stream_internal_oready;
  reg [32-1:0] _stream_conv2d_25_fsm;
  localparam _stream_conv2d_25_fsm_init = 0;
  wire _stream_conv2d_25_run_flag;
  reg _stream_conv2d_25_source_start;
  wire _stream_conv2d_25_source_stop;
  reg _stream_conv2d_25_source_busy;
  wire _stream_conv2d_25_sink_start;
  wire _stream_conv2d_25_sink_stop;
  wire _stream_conv2d_25_sink_busy;
  wire _stream_conv2d_25_busy;
  reg _stream_conv2d_25_busy_reg;
  wire _stream_conv2d_25_is_root;
  assign _stream_conv2d_25_is_root = 1;
  reg [10-1:0] _stream_conv2d_25_parameter_0_next_parameter_data;
  reg [2-1:0] _stream_conv2d_25_parameter_1_next_parameter_data;
  reg [2-1:0] _stream_conv2d_25_parameter_2_next_parameter_data;
  reg [9-1:0] _stream_conv2d_25_parameter_3_next_parameter_data;
  reg [1-1:0] _stream_conv2d_25_parameter_4_next_parameter_data;
  reg [1-1:0] _stream_conv2d_25_parameter_6_next_parameter_data;
  reg _stream_conv2d_25_source_7_idle;
  reg [33-1:0] _stream_conv2d_25_source_7_source_count;
  reg [5-1:0] _stream_conv2d_25_source_7_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_7_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_7_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_7_source_size;
  reg [32-1:0] _stream_conv2d_25_source_7_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_7_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_7_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_7_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_7_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_7_source_ram_raddr;
  reg _stream_conv2d_25_source_7_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_7_source_ram_rdata;
  reg _stream_conv2d_25_source_7_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_7_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_7_source_empty_data;
  reg [1-1:0] _stream_conv2d_25_parameter_8_next_parameter_data;
  reg _stream_conv2d_25_source_9_idle;
  reg [33-1:0] _stream_conv2d_25_source_9_source_count;
  reg [5-1:0] _stream_conv2d_25_source_9_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_9_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_9_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_9_source_size;
  reg [32-1:0] _stream_conv2d_25_source_9_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_9_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_9_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_9_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_9_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_9_source_ram_raddr;
  reg _stream_conv2d_25_source_9_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_9_source_ram_rdata;
  reg _stream_conv2d_25_source_9_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_9_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_9_source_empty_data;
  reg [1-1:0] _stream_conv2d_25_parameter_10_next_parameter_data;
  reg _stream_conv2d_25_source_11_idle;
  reg [33-1:0] _stream_conv2d_25_source_11_source_count;
  reg [5-1:0] _stream_conv2d_25_source_11_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_11_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_11_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_11_source_size;
  reg [32-1:0] _stream_conv2d_25_source_11_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_11_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_11_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_11_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_11_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_11_source_ram_raddr;
  reg _stream_conv2d_25_source_11_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_11_source_ram_rdata;
  reg _stream_conv2d_25_source_11_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_11_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_11_source_empty_data;
  reg [1-1:0] _stream_conv2d_25_parameter_12_next_parameter_data;
  reg _stream_conv2d_25_source_13_idle;
  reg [33-1:0] _stream_conv2d_25_source_13_source_count;
  reg [5-1:0] _stream_conv2d_25_source_13_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_13_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_13_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_13_source_size;
  reg [32-1:0] _stream_conv2d_25_source_13_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_13_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_13_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_13_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_13_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_13_source_ram_raddr;
  reg _stream_conv2d_25_source_13_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_13_source_ram_rdata;
  reg _stream_conv2d_25_source_13_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_13_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_13_source_empty_data;
  reg [1-1:0] _stream_conv2d_25_parameter_14_next_parameter_data;
  reg _stream_conv2d_25_source_15_idle;
  reg [33-1:0] _stream_conv2d_25_source_15_source_count;
  reg [5-1:0] _stream_conv2d_25_source_15_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_15_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_15_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_15_source_size;
  reg [32-1:0] _stream_conv2d_25_source_15_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_15_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_15_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_15_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_15_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_15_source_ram_raddr;
  reg _stream_conv2d_25_source_15_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_15_source_ram_rdata;
  reg _stream_conv2d_25_source_15_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_15_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_15_source_empty_data;
  reg [1-1:0] _stream_conv2d_25_parameter_16_next_parameter_data;
  reg [1-1:0] _stream_conv2d_25_parameter_17_next_parameter_data;
  reg [5-1:0] _stream_conv2d_25_parameter_18_next_parameter_data;
  reg [1-1:0] _stream_conv2d_25_parameter_19_next_parameter_data;
  reg _stream_conv2d_25_source_20_idle;
  reg [33-1:0] _stream_conv2d_25_source_20_source_count;
  reg [5-1:0] _stream_conv2d_25_source_20_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_20_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_20_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_20_source_size;
  reg [32-1:0] _stream_conv2d_25_source_20_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_20_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_20_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_20_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_20_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_20_source_ram_raddr;
  reg _stream_conv2d_25_source_20_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_20_source_ram_rdata;
  reg _stream_conv2d_25_source_20_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_20_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_20_source_empty_data;
  reg _stream_conv2d_25_source_21_idle;
  reg [33-1:0] _stream_conv2d_25_source_21_source_count;
  reg [5-1:0] _stream_conv2d_25_source_21_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_21_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_21_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_21_source_size;
  reg [32-1:0] _stream_conv2d_25_source_21_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_21_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_21_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_21_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_21_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_21_source_ram_raddr;
  reg _stream_conv2d_25_source_21_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_21_source_ram_rdata;
  reg _stream_conv2d_25_source_21_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_21_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_21_source_empty_data;
  reg _stream_conv2d_25_source_22_idle;
  reg [33-1:0] _stream_conv2d_25_source_22_source_count;
  reg [5-1:0] _stream_conv2d_25_source_22_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_22_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_22_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_22_source_size;
  reg [32-1:0] _stream_conv2d_25_source_22_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_22_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_22_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_22_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_22_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_22_source_ram_raddr;
  reg _stream_conv2d_25_source_22_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_22_source_ram_rdata;
  reg _stream_conv2d_25_source_22_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_22_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_22_source_empty_data;
  reg _stream_conv2d_25_source_23_idle;
  reg [33-1:0] _stream_conv2d_25_source_23_source_count;
  reg [5-1:0] _stream_conv2d_25_source_23_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_23_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_23_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_23_source_size;
  reg [32-1:0] _stream_conv2d_25_source_23_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_23_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_23_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_23_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_23_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_23_source_ram_raddr;
  reg _stream_conv2d_25_source_23_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_23_source_ram_rdata;
  reg _stream_conv2d_25_source_23_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_23_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_23_source_empty_data;
  reg _stream_conv2d_25_source_24_idle;
  reg [33-1:0] _stream_conv2d_25_source_24_source_count;
  reg [5-1:0] _stream_conv2d_25_source_24_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_24_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_24_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_24_source_size;
  reg [32-1:0] _stream_conv2d_25_source_24_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_24_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_24_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_24_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_24_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_24_source_ram_raddr;
  reg _stream_conv2d_25_source_24_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_24_source_ram_rdata;
  reg _stream_conv2d_25_source_24_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_24_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_24_source_empty_data;
  reg _stream_conv2d_25_source_25_idle;
  reg [33-1:0] _stream_conv2d_25_source_25_source_count;
  reg [5-1:0] _stream_conv2d_25_source_25_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_25_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_25_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_25_source_size;
  reg [32-1:0] _stream_conv2d_25_source_25_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_25_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_25_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_25_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_25_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_25_source_ram_raddr;
  reg _stream_conv2d_25_source_25_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_25_source_ram_rdata;
  reg _stream_conv2d_25_source_25_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_25_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_25_source_empty_data;
  reg _stream_conv2d_25_source_26_idle;
  reg [33-1:0] _stream_conv2d_25_source_26_source_count;
  reg [5-1:0] _stream_conv2d_25_source_26_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_26_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_26_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_26_source_size;
  reg [32-1:0] _stream_conv2d_25_source_26_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_26_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_26_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_26_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_26_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_26_source_ram_raddr;
  reg _stream_conv2d_25_source_26_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_26_source_ram_rdata;
  reg _stream_conv2d_25_source_26_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_26_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_26_source_empty_data;
  reg _stream_conv2d_25_source_27_idle;
  reg [33-1:0] _stream_conv2d_25_source_27_source_count;
  reg [5-1:0] _stream_conv2d_25_source_27_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_27_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_27_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_27_source_size;
  reg [32-1:0] _stream_conv2d_25_source_27_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_27_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_27_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_27_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_27_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_27_source_ram_raddr;
  reg _stream_conv2d_25_source_27_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_27_source_ram_rdata;
  reg _stream_conv2d_25_source_27_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_27_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_27_source_empty_data;
  reg _stream_conv2d_25_source_28_idle;
  reg [33-1:0] _stream_conv2d_25_source_28_source_count;
  reg [5-1:0] _stream_conv2d_25_source_28_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_28_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_28_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_28_source_size;
  reg [32-1:0] _stream_conv2d_25_source_28_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_28_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_28_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_28_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_28_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_28_source_ram_raddr;
  reg _stream_conv2d_25_source_28_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_28_source_ram_rdata;
  reg _stream_conv2d_25_source_28_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_28_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_28_source_empty_data;
  reg _stream_conv2d_25_source_29_idle;
  reg [33-1:0] _stream_conv2d_25_source_29_source_count;
  reg [5-1:0] _stream_conv2d_25_source_29_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_29_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_29_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_29_source_size;
  reg [32-1:0] _stream_conv2d_25_source_29_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_29_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_29_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_29_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_29_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_29_source_ram_raddr;
  reg _stream_conv2d_25_source_29_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_29_source_ram_rdata;
  reg _stream_conv2d_25_source_29_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_29_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_29_source_empty_data;
  reg _stream_conv2d_25_source_30_idle;
  reg [33-1:0] _stream_conv2d_25_source_30_source_count;
  reg [5-1:0] _stream_conv2d_25_source_30_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_30_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_30_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_30_source_size;
  reg [32-1:0] _stream_conv2d_25_source_30_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_30_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_30_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_30_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_30_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_30_source_ram_raddr;
  reg _stream_conv2d_25_source_30_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_30_source_ram_rdata;
  reg _stream_conv2d_25_source_30_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_30_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_30_source_empty_data;
  reg _stream_conv2d_25_source_31_idle;
  reg [33-1:0] _stream_conv2d_25_source_31_source_count;
  reg [5-1:0] _stream_conv2d_25_source_31_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_31_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_31_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_31_source_size;
  reg [32-1:0] _stream_conv2d_25_source_31_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_31_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_31_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_31_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_31_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_31_source_ram_raddr;
  reg _stream_conv2d_25_source_31_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_31_source_ram_rdata;
  reg _stream_conv2d_25_source_31_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_31_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_31_source_empty_data;
  reg _stream_conv2d_25_source_32_idle;
  reg [33-1:0] _stream_conv2d_25_source_32_source_count;
  reg [5-1:0] _stream_conv2d_25_source_32_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_32_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_32_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_32_source_size;
  reg [32-1:0] _stream_conv2d_25_source_32_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_32_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_32_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_32_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_32_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_32_source_ram_raddr;
  reg _stream_conv2d_25_source_32_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_32_source_ram_rdata;
  reg _stream_conv2d_25_source_32_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_32_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_32_source_empty_data;
  reg _stream_conv2d_25_source_33_idle;
  reg [33-1:0] _stream_conv2d_25_source_33_source_count;
  reg [5-1:0] _stream_conv2d_25_source_33_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_33_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_33_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_33_source_size;
  reg [32-1:0] _stream_conv2d_25_source_33_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_33_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_33_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_33_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_33_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_33_source_ram_raddr;
  reg _stream_conv2d_25_source_33_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_33_source_ram_rdata;
  reg _stream_conv2d_25_source_33_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_33_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_33_source_empty_data;
  reg _stream_conv2d_25_source_34_idle;
  reg [33-1:0] _stream_conv2d_25_source_34_source_count;
  reg [5-1:0] _stream_conv2d_25_source_34_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_34_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_34_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_34_source_size;
  reg [32-1:0] _stream_conv2d_25_source_34_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_34_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_34_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_34_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_34_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_34_source_ram_raddr;
  reg _stream_conv2d_25_source_34_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_34_source_ram_rdata;
  reg _stream_conv2d_25_source_34_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_34_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_34_source_empty_data;
  reg _stream_conv2d_25_source_35_idle;
  reg [33-1:0] _stream_conv2d_25_source_35_source_count;
  reg [5-1:0] _stream_conv2d_25_source_35_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_35_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_35_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_35_source_size;
  reg [32-1:0] _stream_conv2d_25_source_35_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_35_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_35_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_35_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_35_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_35_source_ram_raddr;
  reg _stream_conv2d_25_source_35_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_35_source_ram_rdata;
  reg _stream_conv2d_25_source_35_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_35_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_35_source_empty_data;
  reg _stream_conv2d_25_source_36_idle;
  reg [33-1:0] _stream_conv2d_25_source_36_source_count;
  reg [5-1:0] _stream_conv2d_25_source_36_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_36_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_36_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_36_source_size;
  reg [32-1:0] _stream_conv2d_25_source_36_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_36_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_36_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_36_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_36_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_36_source_ram_raddr;
  reg _stream_conv2d_25_source_36_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_36_source_ram_rdata;
  reg _stream_conv2d_25_source_36_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_36_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_36_source_empty_data;
  reg _stream_conv2d_25_source_37_idle;
  reg [33-1:0] _stream_conv2d_25_source_37_source_count;
  reg [5-1:0] _stream_conv2d_25_source_37_source_mode;
  reg [16-1:0] _stream_conv2d_25_source_37_source_generator_id;
  reg [32-1:0] _stream_conv2d_25_source_37_source_offset;
  reg [33-1:0] _stream_conv2d_25_source_37_source_size;
  reg [32-1:0] _stream_conv2d_25_source_37_source_stride;
  reg [32-1:0] _stream_conv2d_25_source_37_source_offset_buf;
  reg [33-1:0] _stream_conv2d_25_source_37_source_size_buf;
  reg [32-1:0] _stream_conv2d_25_source_37_source_stride_buf;
  reg [8-1:0] _stream_conv2d_25_source_37_source_sel;
  reg [32-1:0] _stream_conv2d_25_source_37_source_ram_raddr;
  reg _stream_conv2d_25_source_37_source_ram_renable;
  wire [32-1:0] _stream_conv2d_25_source_37_source_ram_rdata;
  reg _stream_conv2d_25_source_37_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_25_source_37_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_25_source_37_source_empty_data;
  wire signed [32-1:0] mul_4_x_data;
  wire signed [32-1:0] mul_4_y_data;
  wire [6-1:0] mul_4_rshift_data;
  reg __mul_4_stream_ivalid_1;
  reg __mul_4_stream_ivalid_2;
  reg __mul_4_stream_ivalid_3;
  reg __mul_4_stream_ivalid_4;
  reg __mul_4_stream_ivalid_5;
  reg __mul_4_stream_ivalid_6;
  reg __mul_4_stream_ivalid_7;
  reg __mul_4_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_83;
  reg [6-1:0] _minus_data_85;
  reg [1-1:0] _greatereq_data_96;
  reg signed [32-1:0] __delay_data_658__variable_80;
  reg signed [32-1:0] __delay_data_661__variable_81;
  reg [6-1:0] __delay_data_664__variable_82;
  reg signed [66-1:0] _sll_data_87;
  reg [1-1:0] __delay_data_655_greaterthan_83;
  reg [1-1:0] __delay_data_656_greatereq_96;
  reg signed [32-1:0] __delay_data_659__delay_658__variable_80;
  reg signed [32-1:0] __delay_data_662__delay_661__variable_81;
  reg [6-1:0] __delay_data_665__delay_664__variable_82;
  reg signed [64-1:0] _cond_data_93;
  reg [1-1:0] __delay_data_657__delay_656_greatereq_96;
  reg signed [32-1:0] __delay_data_660__delay_659__delay_658__variable_80;
  reg signed [32-1:0] __delay_data_663__delay_662__delay_661__variable_81;
  reg [6-1:0] __delay_data_666__delay_665__delay_664__variable_82;
  wire signed [32-1:0] _uminus_data_95;
  assign _uminus_data_95 = -_cond_data_93;
  wire signed [32-1:0] _cond_data_98;
  assign _cond_data_98 = (__delay_data_657__delay_656_greatereq_96)? _cond_data_93 : _uminus_data_95;
  wire signed [64-1:0] __muladd_madd_odata_99;
  reg signed [64-1:0] __muladd_madd_odata_reg_99;
  wire signed [64-1:0] __muladd_data_99;
  assign __muladd_data_99 = __muladd_madd_odata_reg_99;
  wire __muladd_madd_update_99;
  assign __muladd_madd_update_99 = _mul_4_stream_oready;

  madd_0
  __muladd_madd_99
  (
    .CLK(CLK),
    .update(__muladd_madd_update_99),
    .a(__delay_data_660__delay_659__delay_658__variable_80),
    .b(__delay_data_663__delay_662__delay_661__variable_81),
    .c(_cond_data_98),
    .d(__muladd_madd_odata_99)
  );

  reg [6-1:0] __delay_data_667__delay_666__delay_665__delay_664__variable_82;
  reg [6-1:0] __delay_data_668__delay_667__delay_666__delay_665____variable_82;
  reg [6-1:0] __delay_data_669__delay_668__delay_667__delay_666____variable_82;
  reg [6-1:0] __delay_data_670__delay_669__delay_668__delay_667____variable_82;
  reg signed [64-1:0] _sra_data_100;
  wire signed [64-1:0] mul_4_z_data;
  assign mul_4_z_data = _sra_data_100;
  wire signed [32-1:0] mul_5_x_data;
  wire signed [32-1:0] mul_5_y_data;
  wire [6-1:0] mul_5_rshift_data;
  reg __mul_5_stream_ivalid_1;
  reg __mul_5_stream_ivalid_2;
  reg __mul_5_stream_ivalid_3;
  reg __mul_5_stream_ivalid_4;
  reg __mul_5_stream_ivalid_5;
  reg __mul_5_stream_ivalid_6;
  reg __mul_5_stream_ivalid_7;
  reg __mul_5_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_104;
  reg [6-1:0] _minus_data_106;
  reg [1-1:0] _greatereq_data_117;
  reg signed [32-1:0] __delay_data_677__variable_101;
  reg signed [32-1:0] __delay_data_680__variable_102;
  reg [6-1:0] __delay_data_683__variable_103;
  reg signed [66-1:0] _sll_data_108;
  reg [1-1:0] __delay_data_674_greaterthan_104;
  reg [1-1:0] __delay_data_675_greatereq_117;
  reg signed [32-1:0] __delay_data_678__delay_677__variable_101;
  reg signed [32-1:0] __delay_data_681__delay_680__variable_102;
  reg [6-1:0] __delay_data_684__delay_683__variable_103;
  reg signed [64-1:0] _cond_data_114;
  reg [1-1:0] __delay_data_676__delay_675_greatereq_117;
  reg signed [32-1:0] __delay_data_679__delay_678__delay_677__variable_101;
  reg signed [32-1:0] __delay_data_682__delay_681__delay_680__variable_102;
  reg [6-1:0] __delay_data_685__delay_684__delay_683__variable_103;
  wire signed [32-1:0] _uminus_data_116;
  assign _uminus_data_116 = -_cond_data_114;
  wire signed [32-1:0] _cond_data_119;
  assign _cond_data_119 = (__delay_data_676__delay_675_greatereq_117)? _cond_data_114 : _uminus_data_116;
  wire signed [64-1:0] __muladd_madd_odata_120;
  reg signed [64-1:0] __muladd_madd_odata_reg_120;
  wire signed [64-1:0] __muladd_data_120;
  assign __muladd_data_120 = __muladd_madd_odata_reg_120;
  wire __muladd_madd_update_120;
  assign __muladd_madd_update_120 = _mul_5_stream_oready;

  madd_1
  __muladd_madd_120
  (
    .CLK(CLK),
    .update(__muladd_madd_update_120),
    .a(__delay_data_679__delay_678__delay_677__variable_101),
    .b(__delay_data_682__delay_681__delay_680__variable_102),
    .c(_cond_data_119),
    .d(__muladd_madd_odata_120)
  );

  reg [6-1:0] __delay_data_686__delay_685__delay_684____variable_103;
  reg [6-1:0] __delay_data_687__delay_686__delay_685____variable_103;
  reg [6-1:0] __delay_data_688__delay_687__delay_686____variable_103;
  reg [6-1:0] __delay_data_689__delay_688__delay_687____variable_103;
  reg signed [64-1:0] _sra_data_121;
  wire signed [64-1:0] mul_5_z_data;
  assign mul_5_z_data = _sra_data_121;
  wire signed [32-1:0] mul_6_x_data;
  wire signed [32-1:0] mul_6_y_data;
  wire [6-1:0] mul_6_rshift_data;
  reg __mul_6_stream_ivalid_1;
  reg __mul_6_stream_ivalid_2;
  reg __mul_6_stream_ivalid_3;
  reg __mul_6_stream_ivalid_4;
  reg __mul_6_stream_ivalid_5;
  reg __mul_6_stream_ivalid_6;
  reg __mul_6_stream_ivalid_7;
  reg __mul_6_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_125;
  reg [6-1:0] _minus_data_127;
  reg [1-1:0] _greatereq_data_138;
  reg signed [32-1:0] __delay_data_696__variable_122;
  reg signed [32-1:0] __delay_data_699__variable_123;
  reg [6-1:0] __delay_data_702__variable_124;
  reg signed [66-1:0] _sll_data_129;
  reg [1-1:0] __delay_data_693_greaterthan_125;
  reg [1-1:0] __delay_data_694_greatereq_138;
  reg signed [32-1:0] __delay_data_697__delay_696__variable_122;
  reg signed [32-1:0] __delay_data_700__delay_699__variable_123;
  reg [6-1:0] __delay_data_703__delay_702__variable_124;
  reg signed [64-1:0] _cond_data_135;
  reg [1-1:0] __delay_data_695__delay_694_greatereq_138;
  reg signed [32-1:0] __delay_data_698__delay_697__delay_696__variable_122;
  reg signed [32-1:0] __delay_data_701__delay_700__delay_699__variable_123;
  reg [6-1:0] __delay_data_704__delay_703__delay_702__variable_124;
  wire signed [32-1:0] _uminus_data_137;
  assign _uminus_data_137 = -_cond_data_135;
  wire signed [32-1:0] _cond_data_140;
  assign _cond_data_140 = (__delay_data_695__delay_694_greatereq_138)? _cond_data_135 : _uminus_data_137;
  wire signed [64-1:0] __muladd_madd_odata_141;
  reg signed [64-1:0] __muladd_madd_odata_reg_141;
  wire signed [64-1:0] __muladd_data_141;
  assign __muladd_data_141 = __muladd_madd_odata_reg_141;
  wire __muladd_madd_update_141;
  assign __muladd_madd_update_141 = _mul_6_stream_oready;

  madd_2
  __muladd_madd_141
  (
    .CLK(CLK),
    .update(__muladd_madd_update_141),
    .a(__delay_data_698__delay_697__delay_696__variable_122),
    .b(__delay_data_701__delay_700__delay_699__variable_123),
    .c(_cond_data_140),
    .d(__muladd_madd_odata_141)
  );

  reg [6-1:0] __delay_data_705__delay_704__delay_703____variable_124;
  reg [6-1:0] __delay_data_706__delay_705__delay_704____variable_124;
  reg [6-1:0] __delay_data_707__delay_706__delay_705____variable_124;
  reg [6-1:0] __delay_data_708__delay_707__delay_706____variable_124;
  reg signed [64-1:0] _sra_data_142;
  wire signed [64-1:0] mul_6_z_data;
  assign mul_6_z_data = _sra_data_142;
  wire signed [32-1:0] mul_7_x_data;
  wire signed [32-1:0] mul_7_y_data;
  wire [6-1:0] mul_7_rshift_data;
  reg __mul_7_stream_ivalid_1;
  reg __mul_7_stream_ivalid_2;
  reg __mul_7_stream_ivalid_3;
  reg __mul_7_stream_ivalid_4;
  reg __mul_7_stream_ivalid_5;
  reg __mul_7_stream_ivalid_6;
  reg __mul_7_stream_ivalid_7;
  reg __mul_7_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_146;
  reg [6-1:0] _minus_data_148;
  reg [1-1:0] _greatereq_data_159;
  reg signed [32-1:0] __delay_data_715__variable_143;
  reg signed [32-1:0] __delay_data_718__variable_144;
  reg [6-1:0] __delay_data_721__variable_145;
  reg signed [66-1:0] _sll_data_150;
  reg [1-1:0] __delay_data_712_greaterthan_146;
  reg [1-1:0] __delay_data_713_greatereq_159;
  reg signed [32-1:0] __delay_data_716__delay_715__variable_143;
  reg signed [32-1:0] __delay_data_719__delay_718__variable_144;
  reg [6-1:0] __delay_data_722__delay_721__variable_145;
  reg signed [64-1:0] _cond_data_156;
  reg [1-1:0] __delay_data_714__delay_713_greatereq_159;
  reg signed [32-1:0] __delay_data_717__delay_716__delay_715__variable_143;
  reg signed [32-1:0] __delay_data_720__delay_719__delay_718__variable_144;
  reg [6-1:0] __delay_data_723__delay_722__delay_721__variable_145;
  wire signed [32-1:0] _uminus_data_158;
  assign _uminus_data_158 = -_cond_data_156;
  wire signed [32-1:0] _cond_data_161;
  assign _cond_data_161 = (__delay_data_714__delay_713_greatereq_159)? _cond_data_156 : _uminus_data_158;
  wire signed [64-1:0] __muladd_madd_odata_162;
  reg signed [64-1:0] __muladd_madd_odata_reg_162;
  wire signed [64-1:0] __muladd_data_162;
  assign __muladd_data_162 = __muladd_madd_odata_reg_162;
  wire __muladd_madd_update_162;
  assign __muladd_madd_update_162 = _mul_7_stream_oready;

  madd_3
  __muladd_madd_162
  (
    .CLK(CLK),
    .update(__muladd_madd_update_162),
    .a(__delay_data_717__delay_716__delay_715__variable_143),
    .b(__delay_data_720__delay_719__delay_718__variable_144),
    .c(_cond_data_161),
    .d(__muladd_madd_odata_162)
  );

  reg [6-1:0] __delay_data_724__delay_723__delay_722____variable_145;
  reg [6-1:0] __delay_data_725__delay_724__delay_723____variable_145;
  reg [6-1:0] __delay_data_726__delay_725__delay_724____variable_145;
  reg [6-1:0] __delay_data_727__delay_726__delay_725____variable_145;
  reg signed [64-1:0] _sra_data_163;
  wire signed [64-1:0] mul_7_z_data;
  assign mul_7_z_data = _sra_data_163;
  wire signed [32-1:0] mul_8_x_data;
  wire signed [32-1:0] mul_8_y_data;
  wire [6-1:0] mul_8_rshift_data;
  reg __mul_8_stream_ivalid_1;
  reg __mul_8_stream_ivalid_2;
  reg __mul_8_stream_ivalid_3;
  reg __mul_8_stream_ivalid_4;
  reg __mul_8_stream_ivalid_5;
  reg __mul_8_stream_ivalid_6;
  reg __mul_8_stream_ivalid_7;
  reg __mul_8_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_167;
  reg [6-1:0] _minus_data_169;
  reg [1-1:0] _greatereq_data_180;
  reg signed [32-1:0] __delay_data_734__variable_164;
  reg signed [32-1:0] __delay_data_737__variable_165;
  reg [6-1:0] __delay_data_740__variable_166;
  reg signed [66-1:0] _sll_data_171;
  reg [1-1:0] __delay_data_731_greaterthan_167;
  reg [1-1:0] __delay_data_732_greatereq_180;
  reg signed [32-1:0] __delay_data_735__delay_734__variable_164;
  reg signed [32-1:0] __delay_data_738__delay_737__variable_165;
  reg [6-1:0] __delay_data_741__delay_740__variable_166;
  reg signed [64-1:0] _cond_data_177;
  reg [1-1:0] __delay_data_733__delay_732_greatereq_180;
  reg signed [32-1:0] __delay_data_736__delay_735__delay_734__variable_164;
  reg signed [32-1:0] __delay_data_739__delay_738__delay_737__variable_165;
  reg [6-1:0] __delay_data_742__delay_741__delay_740__variable_166;
  wire signed [32-1:0] _uminus_data_179;
  assign _uminus_data_179 = -_cond_data_177;
  wire signed [32-1:0] _cond_data_182;
  assign _cond_data_182 = (__delay_data_733__delay_732_greatereq_180)? _cond_data_177 : _uminus_data_179;
  wire signed [64-1:0] __muladd_madd_odata_183;
  reg signed [64-1:0] __muladd_madd_odata_reg_183;
  wire signed [64-1:0] __muladd_data_183;
  assign __muladd_data_183 = __muladd_madd_odata_reg_183;
  wire __muladd_madd_update_183;
  assign __muladd_madd_update_183 = _mul_8_stream_oready;

  madd_4
  __muladd_madd_183
  (
    .CLK(CLK),
    .update(__muladd_madd_update_183),
    .a(__delay_data_736__delay_735__delay_734__variable_164),
    .b(__delay_data_739__delay_738__delay_737__variable_165),
    .c(_cond_data_182),
    .d(__muladd_madd_odata_183)
  );

  reg [6-1:0] __delay_data_743__delay_742__delay_741____variable_166;
  reg [6-1:0] __delay_data_744__delay_743__delay_742____variable_166;
  reg [6-1:0] __delay_data_745__delay_744__delay_743____variable_166;
  reg [6-1:0] __delay_data_746__delay_745__delay_744____variable_166;
  reg signed [64-1:0] _sra_data_184;
  wire signed [64-1:0] mul_8_z_data;
  assign mul_8_z_data = _sra_data_184;
  wire signed [32-1:0] mul_9_x_data;
  wire signed [32-1:0] mul_9_y_data;
  wire [6-1:0] mul_9_rshift_data;
  reg __mul_9_stream_ivalid_1;
  reg __mul_9_stream_ivalid_2;
  reg __mul_9_stream_ivalid_3;
  reg __mul_9_stream_ivalid_4;
  reg __mul_9_stream_ivalid_5;
  reg __mul_9_stream_ivalid_6;
  reg __mul_9_stream_ivalid_7;
  reg __mul_9_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_188;
  reg [6-1:0] _minus_data_190;
  reg [1-1:0] _greatereq_data_201;
  reg signed [32-1:0] __delay_data_753__variable_185;
  reg signed [32-1:0] __delay_data_756__variable_186;
  reg [6-1:0] __delay_data_759__variable_187;
  reg signed [66-1:0] _sll_data_192;
  reg [1-1:0] __delay_data_750_greaterthan_188;
  reg [1-1:0] __delay_data_751_greatereq_201;
  reg signed [32-1:0] __delay_data_754__delay_753__variable_185;
  reg signed [32-1:0] __delay_data_757__delay_756__variable_186;
  reg [6-1:0] __delay_data_760__delay_759__variable_187;
  reg signed [64-1:0] _cond_data_198;
  reg [1-1:0] __delay_data_752__delay_751_greatereq_201;
  reg signed [32-1:0] __delay_data_755__delay_754__delay_753__variable_185;
  reg signed [32-1:0] __delay_data_758__delay_757__delay_756__variable_186;
  reg [6-1:0] __delay_data_761__delay_760__delay_759__variable_187;
  wire signed [32-1:0] _uminus_data_200;
  assign _uminus_data_200 = -_cond_data_198;
  wire signed [32-1:0] _cond_data_203;
  assign _cond_data_203 = (__delay_data_752__delay_751_greatereq_201)? _cond_data_198 : _uminus_data_200;
  wire signed [64-1:0] __muladd_madd_odata_204;
  reg signed [64-1:0] __muladd_madd_odata_reg_204;
  wire signed [64-1:0] __muladd_data_204;
  assign __muladd_data_204 = __muladd_madd_odata_reg_204;
  wire __muladd_madd_update_204;
  assign __muladd_madd_update_204 = _mul_9_stream_oready;

  madd_5
  __muladd_madd_204
  (
    .CLK(CLK),
    .update(__muladd_madd_update_204),
    .a(__delay_data_755__delay_754__delay_753__variable_185),
    .b(__delay_data_758__delay_757__delay_756__variable_186),
    .c(_cond_data_203),
    .d(__muladd_madd_odata_204)
  );

  reg [6-1:0] __delay_data_762__delay_761__delay_760____variable_187;
  reg [6-1:0] __delay_data_763__delay_762__delay_761____variable_187;
  reg [6-1:0] __delay_data_764__delay_763__delay_762____variable_187;
  reg [6-1:0] __delay_data_765__delay_764__delay_763____variable_187;
  reg signed [64-1:0] _sra_data_205;
  wire signed [64-1:0] mul_9_z_data;
  assign mul_9_z_data = _sra_data_205;
  wire signed [32-1:0] mul_10_x_data;
  wire signed [32-1:0] mul_10_y_data;
  wire [6-1:0] mul_10_rshift_data;
  reg __mul_10_stream_ivalid_1;
  reg __mul_10_stream_ivalid_2;
  reg __mul_10_stream_ivalid_3;
  reg __mul_10_stream_ivalid_4;
  reg __mul_10_stream_ivalid_5;
  reg __mul_10_stream_ivalid_6;
  reg __mul_10_stream_ivalid_7;
  reg __mul_10_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_209;
  reg [6-1:0] _minus_data_211;
  reg [1-1:0] _greatereq_data_222;
  reg signed [32-1:0] __delay_data_772__variable_206;
  reg signed [32-1:0] __delay_data_775__variable_207;
  reg [6-1:0] __delay_data_778__variable_208;
  reg signed [66-1:0] _sll_data_213;
  reg [1-1:0] __delay_data_769_greaterthan_209;
  reg [1-1:0] __delay_data_770_greatereq_222;
  reg signed [32-1:0] __delay_data_773__delay_772__variable_206;
  reg signed [32-1:0] __delay_data_776__delay_775__variable_207;
  reg [6-1:0] __delay_data_779__delay_778__variable_208;
  reg signed [64-1:0] _cond_data_219;
  reg [1-1:0] __delay_data_771__delay_770_greatereq_222;
  reg signed [32-1:0] __delay_data_774__delay_773__delay_772__variable_206;
  reg signed [32-1:0] __delay_data_777__delay_776__delay_775__variable_207;
  reg [6-1:0] __delay_data_780__delay_779__delay_778__variable_208;
  wire signed [32-1:0] _uminus_data_221;
  assign _uminus_data_221 = -_cond_data_219;
  wire signed [32-1:0] _cond_data_224;
  assign _cond_data_224 = (__delay_data_771__delay_770_greatereq_222)? _cond_data_219 : _uminus_data_221;
  wire signed [64-1:0] __muladd_madd_odata_225;
  reg signed [64-1:0] __muladd_madd_odata_reg_225;
  wire signed [64-1:0] __muladd_data_225;
  assign __muladd_data_225 = __muladd_madd_odata_reg_225;
  wire __muladd_madd_update_225;
  assign __muladd_madd_update_225 = _mul_10_stream_oready;

  madd_6
  __muladd_madd_225
  (
    .CLK(CLK),
    .update(__muladd_madd_update_225),
    .a(__delay_data_774__delay_773__delay_772__variable_206),
    .b(__delay_data_777__delay_776__delay_775__variable_207),
    .c(_cond_data_224),
    .d(__muladd_madd_odata_225)
  );

  reg [6-1:0] __delay_data_781__delay_780__delay_779____variable_208;
  reg [6-1:0] __delay_data_782__delay_781__delay_780____variable_208;
  reg [6-1:0] __delay_data_783__delay_782__delay_781____variable_208;
  reg [6-1:0] __delay_data_784__delay_783__delay_782____variable_208;
  reg signed [64-1:0] _sra_data_226;
  wire signed [64-1:0] mul_10_z_data;
  assign mul_10_z_data = _sra_data_226;
  wire signed [32-1:0] mul_11_x_data;
  wire signed [32-1:0] mul_11_y_data;
  wire [6-1:0] mul_11_rshift_data;
  reg __mul_11_stream_ivalid_1;
  reg __mul_11_stream_ivalid_2;
  reg __mul_11_stream_ivalid_3;
  reg __mul_11_stream_ivalid_4;
  reg __mul_11_stream_ivalid_5;
  reg __mul_11_stream_ivalid_6;
  reg __mul_11_stream_ivalid_7;
  reg __mul_11_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_230;
  reg [6-1:0] _minus_data_232;
  reg [1-1:0] _greatereq_data_243;
  reg signed [32-1:0] __delay_data_791__variable_227;
  reg signed [32-1:0] __delay_data_794__variable_228;
  reg [6-1:0] __delay_data_797__variable_229;
  reg signed [66-1:0] _sll_data_234;
  reg [1-1:0] __delay_data_788_greaterthan_230;
  reg [1-1:0] __delay_data_789_greatereq_243;
  reg signed [32-1:0] __delay_data_792__delay_791__variable_227;
  reg signed [32-1:0] __delay_data_795__delay_794__variable_228;
  reg [6-1:0] __delay_data_798__delay_797__variable_229;
  reg signed [64-1:0] _cond_data_240;
  reg [1-1:0] __delay_data_790__delay_789_greatereq_243;
  reg signed [32-1:0] __delay_data_793__delay_792__delay_791__variable_227;
  reg signed [32-1:0] __delay_data_796__delay_795__delay_794__variable_228;
  reg [6-1:0] __delay_data_799__delay_798__delay_797__variable_229;
  wire signed [32-1:0] _uminus_data_242;
  assign _uminus_data_242 = -_cond_data_240;
  wire signed [32-1:0] _cond_data_245;
  assign _cond_data_245 = (__delay_data_790__delay_789_greatereq_243)? _cond_data_240 : _uminus_data_242;
  wire signed [64-1:0] __muladd_madd_odata_246;
  reg signed [64-1:0] __muladd_madd_odata_reg_246;
  wire signed [64-1:0] __muladd_data_246;
  assign __muladd_data_246 = __muladd_madd_odata_reg_246;
  wire __muladd_madd_update_246;
  assign __muladd_madd_update_246 = _mul_11_stream_oready;

  madd_7
  __muladd_madd_246
  (
    .CLK(CLK),
    .update(__muladd_madd_update_246),
    .a(__delay_data_793__delay_792__delay_791__variable_227),
    .b(__delay_data_796__delay_795__delay_794__variable_228),
    .c(_cond_data_245),
    .d(__muladd_madd_odata_246)
  );

  reg [6-1:0] __delay_data_800__delay_799__delay_798____variable_229;
  reg [6-1:0] __delay_data_801__delay_800__delay_799____variable_229;
  reg [6-1:0] __delay_data_802__delay_801__delay_800____variable_229;
  reg [6-1:0] __delay_data_803__delay_802__delay_801____variable_229;
  reg signed [64-1:0] _sra_data_247;
  wire signed [64-1:0] mul_11_z_data;
  assign mul_11_z_data = _sra_data_247;
  wire signed [32-1:0] mul_12_x_data;
  wire signed [32-1:0] mul_12_y_data;
  wire [6-1:0] mul_12_rshift_data;
  reg __mul_12_stream_ivalid_1;
  reg __mul_12_stream_ivalid_2;
  reg __mul_12_stream_ivalid_3;
  reg __mul_12_stream_ivalid_4;
  reg __mul_12_stream_ivalid_5;
  reg __mul_12_stream_ivalid_6;
  reg __mul_12_stream_ivalid_7;
  reg __mul_12_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_251;
  reg [6-1:0] _minus_data_253;
  reg [1-1:0] _greatereq_data_264;
  reg signed [32-1:0] __delay_data_810__variable_248;
  reg signed [32-1:0] __delay_data_813__variable_249;
  reg [6-1:0] __delay_data_816__variable_250;
  reg signed [66-1:0] _sll_data_255;
  reg [1-1:0] __delay_data_807_greaterthan_251;
  reg [1-1:0] __delay_data_808_greatereq_264;
  reg signed [32-1:0] __delay_data_811__delay_810__variable_248;
  reg signed [32-1:0] __delay_data_814__delay_813__variable_249;
  reg [6-1:0] __delay_data_817__delay_816__variable_250;
  reg signed [64-1:0] _cond_data_261;
  reg [1-1:0] __delay_data_809__delay_808_greatereq_264;
  reg signed [32-1:0] __delay_data_812__delay_811__delay_810__variable_248;
  reg signed [32-1:0] __delay_data_815__delay_814__delay_813__variable_249;
  reg [6-1:0] __delay_data_818__delay_817__delay_816__variable_250;
  wire signed [32-1:0] _uminus_data_263;
  assign _uminus_data_263 = -_cond_data_261;
  wire signed [32-1:0] _cond_data_266;
  assign _cond_data_266 = (__delay_data_809__delay_808_greatereq_264)? _cond_data_261 : _uminus_data_263;
  wire signed [64-1:0] __muladd_madd_odata_267;
  reg signed [64-1:0] __muladd_madd_odata_reg_267;
  wire signed [64-1:0] __muladd_data_267;
  assign __muladd_data_267 = __muladd_madd_odata_reg_267;
  wire __muladd_madd_update_267;
  assign __muladd_madd_update_267 = _mul_12_stream_oready;

  madd_8
  __muladd_madd_267
  (
    .CLK(CLK),
    .update(__muladd_madd_update_267),
    .a(__delay_data_812__delay_811__delay_810__variable_248),
    .b(__delay_data_815__delay_814__delay_813__variable_249),
    .c(_cond_data_266),
    .d(__muladd_madd_odata_267)
  );

  reg [6-1:0] __delay_data_819__delay_818__delay_817____variable_250;
  reg [6-1:0] __delay_data_820__delay_819__delay_818____variable_250;
  reg [6-1:0] __delay_data_821__delay_820__delay_819____variable_250;
  reg [6-1:0] __delay_data_822__delay_821__delay_820____variable_250;
  reg signed [64-1:0] _sra_data_268;
  wire signed [64-1:0] mul_12_z_data;
  assign mul_12_z_data = _sra_data_268;
  wire signed [128-1:0] add_tree_2_var0_data;
  wire signed [128-1:0] add_tree_2_var1_data;
  wire signed [128-1:0] add_tree_2_var2_data;
  wire signed [128-1:0] add_tree_2_var3_data;
  wire signed [128-1:0] add_tree_2_var4_data;
  wire signed [128-1:0] add_tree_2_var5_data;
  wire signed [128-1:0] add_tree_2_var6_data;
  wire signed [128-1:0] add_tree_2_var7_data;
  wire signed [128-1:0] add_tree_2_var8_data;
  reg __add_tree_2_stream_ivalid_1;
  reg __add_tree_2_stream_ivalid_2;
  reg signed [128-1:0] __plusn_data_42;
  reg signed [128-1:0] __plusn_data_43;
  reg signed [128-1:0] __plusn_data_44;
  reg signed [128-1:0] __plusn_data_45;
  wire signed [128-1:0] add_tree_2_sum_data;
  assign add_tree_2_sum_data = __plusn_data_45;
  wire signed [128-1:0] acc_1_x_data;
  wire [8-1:0] acc_1_rshift_data;
  wire [32-1:0] acc_1_size_data;
  wire [1-1:0] acc_1__reduce_reset_data;
  reg __acc_1_stream_ivalid_1;
  reg __acc_1_stream_ivalid_2;
  reg __acc_1_stream_ivalid_3;
  reg __acc_1_stream_ivalid_4;
  reg __acc_1_stream_ivalid_5;
  reg [1-1:0] _greaterthan_data_13;
  reg [8-1:0] _minus_data_15;
  reg signed [128-1:0] _reduceadd_data_26;
  reg [33-1:0] _reduceadd_count_26;
  reg _reduceadd_prev_count_max_26;
  wire _reduceadd_reset_cond_26;
  assign _reduceadd_reset_cond_26 = acc_1__reduce_reset_data || _reduceadd_prev_count_max_26;
  wire [33-1:0] _reduceadd_current_count_26;
  assign _reduceadd_current_count_26 = (_reduceadd_reset_cond_26)? 0 : _reduceadd_count_26;
  wire signed [128-1:0] _reduceadd_current_data_26;
  assign _reduceadd_current_data_26 = (_reduceadd_reset_cond_26)? 1'sd0 : _reduceadd_data_26;
  reg [1-1:0] _pulse_data_28;
  reg [33-1:0] _pulse_count_28;
  reg _pulse_prev_count_max_28;
  wire _pulse_reset_cond_28;
  assign _pulse_reset_cond_28 = acc_1__reduce_reset_data || _pulse_prev_count_max_28;
  wire [33-1:0] _pulse_current_count_28;
  assign _pulse_current_count_28 = (_pulse_reset_cond_28)? 0 : _pulse_count_28;
  wire [1-1:0] _pulse_current_data_28;
  assign _pulse_current_data_28 = (_pulse_reset_cond_28)? 1'sd0 : _pulse_data_28;
  reg [8-1:0] __delay_data_831__variable_11;
  reg signed [258-1:0] _sll_data_17;
  reg [1-1:0] __delay_data_828_greaterthan_13;
  reg signed [128-1:0] __delay_data_829_reduceadd_26;
  reg [8-1:0] __delay_data_832__delay_831__variable_11;
  reg [1-1:0] __delay_data_835_pulse_28;
  reg signed [128-1:0] _cond_data_23;
  reg signed [128-1:0] __delay_data_830__delay_829_reduceadd_26;
  reg [8-1:0] __delay_data_833__delay_832__delay_831__variable_11;
  reg [1-1:0] __delay_data_836__delay_835_pulse_28;
  reg signed [128-1:0] _plus_data_30;
  reg [8-1:0] __delay_data_834__delay_833__delay_832__delay_831__variable_11;
  reg [1-1:0] __delay_data_837__delay_836__delay_835_pulse_28;
  reg signed [128-1:0] _sra_data_31;
  reg [1-1:0] __delay_data_838__delay_837__delay_836__delay_835_pulse_28;
  wire signed [128-1:0] acc_1_sum_data;
  assign acc_1_sum_data = _sra_data_31;
  wire [1-1:0] acc_1_valid_data;
  assign acc_1_valid_data = __delay_data_838__delay_837__delay_836__delay_835_pulse_28;
  wire signed [128-1:0] mul_rshift_round_clip_3_x_data;
  wire signed [32-1:0] mul_rshift_round_clip_3_y_data;
  wire [8-1:0] mul_rshift_round_clip_3_rshift_data;
  reg __mul_rshift_round_clip_3_stream_ivalid_1;
  reg __mul_rshift_round_clip_3_stream_ivalid_2;
  reg __mul_rshift_round_clip_3_stream_ivalid_3;
  reg __mul_rshift_round_clip_3_stream_ivalid_4;
  reg __mul_rshift_round_clip_3_stream_ivalid_5;
  reg __mul_rshift_round_clip_3_stream_ivalid_6;
  reg __mul_rshift_round_clip_3_stream_ivalid_7;
  reg __mul_rshift_round_clip_3_stream_ivalid_8;
  wire signed [160-1:0] _times_mul_odata_49;
  reg signed [160-1:0] _times_mul_odata_reg_49;
  wire signed [160-1:0] _times_data_49;
  assign _times_data_49 = _times_mul_odata_reg_49;
  wire _times_mul_update_49;
  assign _times_mul_update_49 = _mul_rshift_round_clip_3_stream_oready;

  multiplier_0
  _times_mul_49
  (
    .CLK(CLK),
    .update(_times_mul_update_49),
    .a(mul_rshift_round_clip_3_x_data),
    .b(mul_rshift_round_clip_3_y_data),
    .c(_times_mul_odata_49)
  );

  wire [8-1:0] _minus_data_52;
  assign _minus_data_52 = mul_rshift_round_clip_3_rshift_data - 2'sd1;
  wire signed [258-1:0] _sll_data_55;
  assign _sll_data_55 = 2'sd1 << _minus_data_52;
  wire [1-1:0] _eq_data_67;
  assign _eq_data_67 = mul_rshift_round_clip_3_rshift_data == 1'sd0;
  reg signed [258-1:0] __delay_data_844_sll_55;
  reg [8-1:0] __delay_data_848__variable_48;
  reg [1-1:0] __delay_data_852_eq_67;
  reg signed [258-1:0] __delay_data_845__delay_844_sll_55;
  reg [8-1:0] __delay_data_849__delay_848__variable_48;
  reg [1-1:0] __delay_data_853__delay_852_eq_67;
  reg signed [258-1:0] __delay_data_846__delay_845__delay_844_sll_55;
  reg [8-1:0] __delay_data_850__delay_849__delay_848__variable_48;
  reg [1-1:0] __delay_data_854__delay_853__delay_852_eq_67;
  reg signed [258-1:0] __delay_data_847__delay_846__delay_845__delay_844_sll_55;
  reg [8-1:0] __delay_data_851__delay_850__delay_849__delay_848__variable_48;
  reg [1-1:0] __delay_data_855__delay_854__delay_853__delay_852_eq_67;
  wire [1-1:0] _pointer_data_50;
  assign _pointer_data_50 = _times_data_49[9'sd159];
  wire signed [2-1:0] _cond_data_62;
  assign _cond_data_62 = (_pointer_data_50)? -2'sd1 : 1'sd0;
  wire signed [161-1:0] _plus_data_63;
  assign _plus_data_63 = _times_data_49 + __delay_data_847__delay_846__delay_845__delay_844_sll_55;
  wire signed [161-1:0] _plus_data_64;
  assign _plus_data_64 = _plus_data_63 + _cond_data_62;
  wire signed [160-1:0] _sra_data_65;
  assign _sra_data_65 = _plus_data_64 >>> __delay_data_851__delay_850__delay_849__delay_848__variable_48;
  reg signed [160-1:0] _cond_data_68;
  reg [1-1:0] _greaterthan_data_69;
  reg [1-1:0] _lessthan_data_73;
  reg [1-1:0] _greatereq_data_77;
  reg signed [160-1:0] __delay_data_856_cond_68;
  reg signed [160-1:0] _cond_data_71;
  reg signed [160-1:0] _cond_data_75;
  reg [1-1:0] __delay_data_857_greatereq_77;
  reg signed [32-1:0] _cond_data_79;
  wire signed [32-1:0] mul_rshift_round_clip_3_z_data;
  assign mul_rshift_round_clip_3_z_data = _cond_data_79;
  reg [33-1:0] _stream_conv2d_25_sink_50_sink_count;
  reg [5-1:0] _stream_conv2d_25_sink_50_sink_mode;
  reg [16-1:0] _stream_conv2d_25_sink_50_sink_generator_id;
  reg [32-1:0] _stream_conv2d_25_sink_50_sink_offset;
  reg [33-1:0] _stream_conv2d_25_sink_50_sink_size;
  reg [32-1:0] _stream_conv2d_25_sink_50_sink_stride;
  reg [32-1:0] _stream_conv2d_25_sink_50_sink_offset_buf;
  reg [33-1:0] _stream_conv2d_25_sink_50_sink_size_buf;
  reg [32-1:0] _stream_conv2d_25_sink_50_sink_stride_buf;
  reg [8-1:0] _stream_conv2d_25_sink_50_sink_sel;
  reg [32-1:0] _stream_conv2d_25_sink_50_sink_waddr;
  reg _stream_conv2d_25_sink_50_sink_wenable;
  reg [32-1:0] _stream_conv2d_25_sink_50_sink_wdata;
  reg _stream_conv2d_25_sink_50_sink_fifo_enq;
  reg [32-1:0] _stream_conv2d_25_sink_50_sink_fifo_wdata;
  reg [32-1:0] _stream_conv2d_25_sink_50_sink_immediate;
  reg [33-1:0] _stream_conv2d_25_sink_51_sink_count;
  reg [5-1:0] _stream_conv2d_25_sink_51_sink_mode;
  reg [16-1:0] _stream_conv2d_25_sink_51_sink_generator_id;
  reg [32-1:0] _stream_conv2d_25_sink_51_sink_offset;
  reg [33-1:0] _stream_conv2d_25_sink_51_sink_size;
  reg [32-1:0] _stream_conv2d_25_sink_51_sink_stride;
  reg [32-1:0] _stream_conv2d_25_sink_51_sink_offset_buf;
  reg [33-1:0] _stream_conv2d_25_sink_51_sink_size_buf;
  reg [32-1:0] _stream_conv2d_25_sink_51_sink_stride_buf;
  reg [8-1:0] _stream_conv2d_25_sink_51_sink_sel;
  reg [32-1:0] _stream_conv2d_25_sink_51_sink_waddr;
  reg _stream_conv2d_25_sink_51_sink_wenable;
  reg [1-1:0] _stream_conv2d_25_sink_51_sink_wdata;
  reg _stream_conv2d_25_sink_51_sink_fifo_enq;
  reg [1-1:0] _stream_conv2d_25_sink_51_sink_fifo_wdata;
  reg [1-1:0] _stream_conv2d_25_sink_51_sink_immediate;
  reg _stream_max_pool_serial_27_stream_ivalid;
  wire _stream_max_pool_serial_27_stream_oready;
  wire _stream_max_pool_serial_27_stream_internal_oready;
  assign _stream_max_pool_serial_27_stream_oready = _stream_max_pool_serial_27_stream_internal_oready;
  reg [32-1:0] _stream_max_pool_serial_27_fsm;
  localparam _stream_max_pool_serial_27_fsm_init = 0;
  wire _stream_max_pool_serial_27_run_flag;
  reg _stream_max_pool_serial_27_source_start;
  wire _stream_max_pool_serial_27_source_stop;
  reg _stream_max_pool_serial_27_source_busy;
  wire _stream_max_pool_serial_27_sink_start;
  wire _stream_max_pool_serial_27_sink_stop;
  wire _stream_max_pool_serial_27_sink_busy;
  wire _stream_max_pool_serial_27_busy;
  reg _stream_max_pool_serial_27_busy_reg;
  wire _stream_max_pool_serial_27_is_root;
  assign _stream_max_pool_serial_27_is_root = 1;
  reg [3-1:0] _stream_max_pool_serial_27_parameter_0_next_parameter_data;
  reg _stream_max_pool_serial_27_source_1_idle;
  reg [33-1:0] _stream_max_pool_serial_27_source_1_source_count;
  reg [5-1:0] _stream_max_pool_serial_27_source_1_source_mode;
  reg [16-1:0] _stream_max_pool_serial_27_source_1_source_generator_id;
  reg [32-1:0] _stream_max_pool_serial_27_source_1_source_offset;
  reg [33-1:0] _stream_max_pool_serial_27_source_1_source_size;
  reg [32-1:0] _stream_max_pool_serial_27_source_1_source_stride;
  reg [32-1:0] _stream_max_pool_serial_27_source_1_source_offset_buf;
  reg [33-1:0] _stream_max_pool_serial_27_source_1_source_size_buf;
  reg [32-1:0] _stream_max_pool_serial_27_source_1_source_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_27_source_1_source_sel;
  reg [32-1:0] _stream_max_pool_serial_27_source_1_source_ram_raddr;
  reg _stream_max_pool_serial_27_source_1_source_ram_renable;
  wire [32-1:0] _stream_max_pool_serial_27_source_1_source_ram_rdata;
  reg _stream_max_pool_serial_27_source_1_source_fifo_deq;
  wire [32-1:0] _stream_max_pool_serial_27_source_1_source_fifo_rdata;
  reg [32-1:0] _stream_max_pool_serial_27_source_1_source_empty_data;
  reg [4-1:0] _stream_max_pool_serial_27_parameter_2_next_parameter_data;
  wire signed [32-1:0] _reduce_max_13_x_data;
  wire [32-1:0] _reduce_max_13_size_data;
  wire [1-1:0] _reduce_max_13__reduce_reset_data;
  reg ___reduce_max_13_stream_ivalid_1;
  reg signed [32-1:0] _reducemax_data_272;
  reg [33-1:0] _reducemax_count_272;
  reg _reducemax_prev_count_max_272;
  wire _reducemax_reset_cond_272;
  assign _reducemax_reset_cond_272 = _reduce_max_13__reduce_reset_data || _reducemax_prev_count_max_272;
  wire [33-1:0] _reducemax_current_count_272;
  assign _reducemax_current_count_272 = (_reducemax_reset_cond_272)? 0 : _reducemax_count_272;
  wire signed [32-1:0] _reducemax_current_data_272;
  assign _reducemax_current_data_272 = (_reducemax_reset_cond_272)? -33'sd2147483648 : _reducemax_data_272;
  reg [1-1:0] _pulse_data_274;
  reg [33-1:0] _pulse_count_274;
  reg _pulse_prev_count_max_274;
  wire _pulse_reset_cond_274;
  assign _pulse_reset_cond_274 = _reduce_max_13__reduce_reset_data || _pulse_prev_count_max_274;
  wire [33-1:0] _pulse_current_count_274;
  assign _pulse_current_count_274 = (_pulse_reset_cond_274)? 0 : _pulse_count_274;
  wire [1-1:0] _pulse_current_data_274;
  assign _pulse_current_data_274 = (_pulse_reset_cond_274)? 1'sd0 : _pulse_data_274;
  wire signed [32-1:0] _reduce_max_13_data_data;
  assign _reduce_max_13_data_data = _reducemax_data_272;
  wire [1-1:0] _reduce_max_13_valid_data;
  assign _reduce_max_13_valid_data = _pulse_data_274;
  reg [33-1:0] _stream_max_pool_serial_27_sink_5_sink_count;
  reg [5-1:0] _stream_max_pool_serial_27_sink_5_sink_mode;
  reg [16-1:0] _stream_max_pool_serial_27_sink_5_sink_generator_id;
  reg [32-1:0] _stream_max_pool_serial_27_sink_5_sink_offset;
  reg [33-1:0] _stream_max_pool_serial_27_sink_5_sink_size;
  reg [32-1:0] _stream_max_pool_serial_27_sink_5_sink_stride;
  reg [32-1:0] _stream_max_pool_serial_27_sink_5_sink_offset_buf;
  reg [33-1:0] _stream_max_pool_serial_27_sink_5_sink_size_buf;
  reg [32-1:0] _stream_max_pool_serial_27_sink_5_sink_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_27_sink_5_sink_sel;
  reg [32-1:0] _stream_max_pool_serial_27_sink_5_sink_waddr;
  reg _stream_max_pool_serial_27_sink_5_sink_wenable;
  reg [32-1:0] _stream_max_pool_serial_27_sink_5_sink_wdata;
  reg _stream_max_pool_serial_27_sink_5_sink_fifo_enq;
  reg [32-1:0] _stream_max_pool_serial_27_sink_5_sink_fifo_wdata;
  reg [32-1:0] _stream_max_pool_serial_27_sink_5_sink_immediate;
  reg [33-1:0] _stream_max_pool_serial_27_sink_6_sink_count;
  reg [5-1:0] _stream_max_pool_serial_27_sink_6_sink_mode;
  reg [16-1:0] _stream_max_pool_serial_27_sink_6_sink_generator_id;
  reg [32-1:0] _stream_max_pool_serial_27_sink_6_sink_offset;
  reg [33-1:0] _stream_max_pool_serial_27_sink_6_sink_size;
  reg [32-1:0] _stream_max_pool_serial_27_sink_6_sink_stride;
  reg [32-1:0] _stream_max_pool_serial_27_sink_6_sink_offset_buf;
  reg [33-1:0] _stream_max_pool_serial_27_sink_6_sink_size_buf;
  reg [32-1:0] _stream_max_pool_serial_27_sink_6_sink_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_27_sink_6_sink_sel;
  reg [32-1:0] _stream_max_pool_serial_27_sink_6_sink_waddr;
  reg _stream_max_pool_serial_27_sink_6_sink_wenable;
  reg [1-1:0] _stream_max_pool_serial_27_sink_6_sink_wdata;
  reg _stream_max_pool_serial_27_sink_6_sink_fifo_enq;
  reg [1-1:0] _stream_max_pool_serial_27_sink_6_sink_fifo_wdata;
  reg [1-1:0] _stream_max_pool_serial_27_sink_6_sink_immediate;
  reg _stream_max_pool_47_stream_ivalid;
  wire _stream_max_pool_47_stream_oready;
  wire _stream_max_pool_47_stream_internal_oready;
  assign _stream_max_pool_47_stream_oready = _stream_max_pool_47_stream_internal_oready;
  reg [32-1:0] _stream_max_pool_47_fsm;
  localparam _stream_max_pool_47_fsm_init = 0;
  wire _stream_max_pool_47_run_flag;
  reg _stream_max_pool_47_source_start;
  wire _stream_max_pool_47_source_stop;
  reg _stream_max_pool_47_source_busy;
  wire _stream_max_pool_47_sink_start;
  wire _stream_max_pool_47_sink_stop;
  wire _stream_max_pool_47_sink_busy;
  wire _stream_max_pool_47_busy;
  reg _stream_max_pool_47_busy_reg;
  wire _stream_max_pool_47_is_root;
  assign _stream_max_pool_47_is_root = 1;
  reg [4-1:0] _stream_max_pool_47_parameter_0_next_parameter_data;
  reg _stream_max_pool_47_source_1_idle;
  reg [33-1:0] _stream_max_pool_47_source_1_source_count;
  reg [5-1:0] _stream_max_pool_47_source_1_source_mode;
  reg [16-1:0] _stream_max_pool_47_source_1_source_generator_id;
  reg [32-1:0] _stream_max_pool_47_source_1_source_offset;
  reg [33-1:0] _stream_max_pool_47_source_1_source_size;
  reg [32-1:0] _stream_max_pool_47_source_1_source_stride;
  reg [32-1:0] _stream_max_pool_47_source_1_source_offset_buf;
  reg [33-1:0] _stream_max_pool_47_source_1_source_size_buf;
  reg [32-1:0] _stream_max_pool_47_source_1_source_stride_buf;
  reg [8-1:0] _stream_max_pool_47_source_1_source_sel;
  reg [32-1:0] _stream_max_pool_47_source_1_source_ram_raddr;
  reg _stream_max_pool_47_source_1_source_ram_renable;
  wire [32-1:0] _stream_max_pool_47_source_1_source_ram_rdata;
  reg _stream_max_pool_47_source_1_source_fifo_deq;
  wire [32-1:0] _stream_max_pool_47_source_1_source_fifo_rdata;
  reg [32-1:0] _stream_max_pool_47_source_1_source_empty_data;
  reg _stream_max_pool_47_source_2_idle;
  reg [33-1:0] _stream_max_pool_47_source_2_source_count;
  reg [5-1:0] _stream_max_pool_47_source_2_source_mode;
  reg [16-1:0] _stream_max_pool_47_source_2_source_generator_id;
  reg [32-1:0] _stream_max_pool_47_source_2_source_offset;
  reg [33-1:0] _stream_max_pool_47_source_2_source_size;
  reg [32-1:0] _stream_max_pool_47_source_2_source_stride;
  reg [32-1:0] _stream_max_pool_47_source_2_source_offset_buf;
  reg [33-1:0] _stream_max_pool_47_source_2_source_size_buf;
  reg [32-1:0] _stream_max_pool_47_source_2_source_stride_buf;
  reg [8-1:0] _stream_max_pool_47_source_2_source_sel;
  reg [32-1:0] _stream_max_pool_47_source_2_source_ram_raddr;
  reg _stream_max_pool_47_source_2_source_ram_renable;
  wire [32-1:0] _stream_max_pool_47_source_2_source_ram_rdata;
  reg _stream_max_pool_47_source_2_source_fifo_deq;
  wire [32-1:0] _stream_max_pool_47_source_2_source_fifo_rdata;
  reg [32-1:0] _stream_max_pool_47_source_2_source_empty_data;
  reg _stream_max_pool_47_source_3_idle;
  reg [33-1:0] _stream_max_pool_47_source_3_source_count;
  reg [5-1:0] _stream_max_pool_47_source_3_source_mode;
  reg [16-1:0] _stream_max_pool_47_source_3_source_generator_id;
  reg [32-1:0] _stream_max_pool_47_source_3_source_offset;
  reg [33-1:0] _stream_max_pool_47_source_3_source_size;
  reg [32-1:0] _stream_max_pool_47_source_3_source_stride;
  reg [32-1:0] _stream_max_pool_47_source_3_source_offset_buf;
  reg [33-1:0] _stream_max_pool_47_source_3_source_size_buf;
  reg [32-1:0] _stream_max_pool_47_source_3_source_stride_buf;
  reg [8-1:0] _stream_max_pool_47_source_3_source_sel;
  reg [32-1:0] _stream_max_pool_47_source_3_source_ram_raddr;
  reg _stream_max_pool_47_source_3_source_ram_renable;
  wire [32-1:0] _stream_max_pool_47_source_3_source_ram_rdata;
  reg _stream_max_pool_47_source_3_source_fifo_deq;
  wire [32-1:0] _stream_max_pool_47_source_3_source_fifo_rdata;
  reg [32-1:0] _stream_max_pool_47_source_3_source_empty_data;
  reg _stream_max_pool_47_source_4_idle;
  reg [33-1:0] _stream_max_pool_47_source_4_source_count;
  reg [5-1:0] _stream_max_pool_47_source_4_source_mode;
  reg [16-1:0] _stream_max_pool_47_source_4_source_generator_id;
  reg [32-1:0] _stream_max_pool_47_source_4_source_offset;
  reg [33-1:0] _stream_max_pool_47_source_4_source_size;
  reg [32-1:0] _stream_max_pool_47_source_4_source_stride;
  reg [32-1:0] _stream_max_pool_47_source_4_source_offset_buf;
  reg [33-1:0] _stream_max_pool_47_source_4_source_size_buf;
  reg [32-1:0] _stream_max_pool_47_source_4_source_stride_buf;
  reg [8-1:0] _stream_max_pool_47_source_4_source_sel;
  reg [32-1:0] _stream_max_pool_47_source_4_source_ram_raddr;
  reg _stream_max_pool_47_source_4_source_ram_renable;
  wire [32-1:0] _stream_max_pool_47_source_4_source_ram_rdata;
  reg _stream_max_pool_47_source_4_source_fifo_deq;
  wire [32-1:0] _stream_max_pool_47_source_4_source_fifo_rdata;
  reg [32-1:0] _stream_max_pool_47_source_4_source_empty_data;
  wire signed [32-1:0] _max_0_var0_data;
  wire signed [32-1:0] _max_0_var1_data;
  wire signed [32-1:0] _max_0_var2_data;
  wire signed [32-1:0] _max_0_var3_data;
  reg ___max_0_stream_ivalid_1;
  reg ___max_0_stream_ivalid_2;
  reg ___max_0_stream_ivalid_3;
  reg ___max_0_stream_ivalid_4;
  reg [1-1:0] _greaterthan_data_4;
  reg [1-1:0] _greaterthan_data_6;
  reg signed [32-1:0] __delay_data_938__variable_0;
  reg signed [32-1:0] __delay_data_939__variable_1;
  reg signed [32-1:0] __delay_data_940__variable_2;
  reg signed [32-1:0] __delay_data_941__variable_3;
  reg signed [32-1:0] _cond_data_5;
  reg signed [32-1:0] _cond_data_7;
  reg [1-1:0] _greaterthan_data_8;
  reg signed [32-1:0] __delay_data_942_cond_5;
  reg signed [32-1:0] __delay_data_943_cond_7;
  reg signed [32-1:0] _cond_data_9;
  wire signed [32-1:0] _max_0_val_data;
  assign _max_0_val_data = _cond_data_9;
  reg [33-1:0] _stream_max_pool_47_sink_6_sink_count;
  reg [5-1:0] _stream_max_pool_47_sink_6_sink_mode;
  reg [16-1:0] _stream_max_pool_47_sink_6_sink_generator_id;
  reg [32-1:0] _stream_max_pool_47_sink_6_sink_offset;
  reg [33-1:0] _stream_max_pool_47_sink_6_sink_size;
  reg [32-1:0] _stream_max_pool_47_sink_6_sink_stride;
  reg [32-1:0] _stream_max_pool_47_sink_6_sink_offset_buf;
  reg [33-1:0] _stream_max_pool_47_sink_6_sink_size_buf;
  reg [32-1:0] _stream_max_pool_47_sink_6_sink_stride_buf;
  reg [8-1:0] _stream_max_pool_47_sink_6_sink_sel;
  reg [32-1:0] _stream_max_pool_47_sink_6_sink_waddr;
  reg _stream_max_pool_47_sink_6_sink_wenable;
  reg [32-1:0] _stream_max_pool_47_sink_6_sink_wdata;
  reg _stream_max_pool_47_sink_6_sink_fifo_enq;
  reg [32-1:0] _stream_max_pool_47_sink_6_sink_fifo_wdata;
  reg [32-1:0] _stream_max_pool_47_sink_6_sink_immediate;
  reg [32-1:0] main_fsm;
  localparam main_fsm_init = 0;
  reg [32-1:0] internal_state_counter;
  reg [32-1:0] conv2d_25_objaddr;
  reg [32-1:0] conv2d_25_arg_objaddr_0;
  reg [32-1:0] conv2d_25_arg_objaddr_1;
  reg [32-1:0] conv2d_25_arg_objaddr_2;
  reg [32-1:0] conv2d_25_arg_objaddr_3;
  reg [32-1:0] control_conv2d_25;
  localparam control_conv2d_25_init = 0;
  reg _control_conv2d_25_called;
  wire signed [32-1:0] conv2d_25_act_base_offset;
  reg signed [32-1:0] conv2d_25_act_base_offset_row;
  reg signed [32-1:0] conv2d_25_act_base_offset_bat;
  assign conv2d_25_act_base_offset = conv2d_25_act_base_offset_row + conv2d_25_act_base_offset_bat;
  reg signed [32-1:0] conv2d_25_filter_base_offset;
  reg [32-1:0] conv2d_25_next_stream_num_ops;
  wire signed [32-1:0] conv2d_25_out_base_offset;
  reg signed [32-1:0] conv2d_25_out_base_offset_val;
  reg signed [32-1:0] conv2d_25_out_base_offset_col;
  reg signed [32-1:0] conv2d_25_out_base_offset_row;
  reg signed [32-1:0] conv2d_25_out_base_offset_bat;
  reg signed [32-1:0] conv2d_25_out_base_offset_och;
  assign conv2d_25_out_base_offset = conv2d_25_out_base_offset_val + conv2d_25_out_base_offset_col + conv2d_25_out_base_offset_row + conv2d_25_out_base_offset_bat + conv2d_25_out_base_offset_och;
  reg conv2d_25_dma_flag_0;
  reg conv2d_25_dma_flag_1;
  reg conv2d_25_dma_flag_2;
  reg [32-1:0] conv2d_25_sync_comp_count;
  reg [32-1:0] conv2d_25_sync_out_count;
  reg [32-1:0] conv2d_25_write_count;
  reg [32-1:0] conv2d_25_next_out_write_size;
  reg [32-1:0] conv2d_25_col_count;
  reg [32-1:0] conv2d_25_row_count;
  reg [32-1:0] conv2d_25_bat_count;
  reg [32-1:0] conv2d_25_och_count;
  reg [2-1:0] conv2d_25_col_select;
  reg [2-1:0] conv2d_25_row_select;
  reg [32-1:0] conv2d_25_out_col_count;
  reg [32-1:0] conv2d_25_out_row_count;
  reg [32-1:0] conv2d_25_out_ram_select;
  reg [32-1:0] conv2d_25_prev_col_count;
  reg [32-1:0] conv2d_25_prev_row_count;
  reg [32-1:0] conv2d_25_prev_bat_count;
  reg [32-1:0] conv2d_25_prev_och_count;
  reg [2-1:0] conv2d_25_prev_row_select;
  reg [32-1:0] conv2d_25_stream_act_local_0;
  reg [32-1:0] conv2d_25_stream_act_local_1;
  reg [32-1:0] conv2d_25_stream_act_local_2;
  reg [32-1:0] conv2d_25_stream_act_local_3;
  reg [32-1:0] conv2d_25_stream_act_local_4;
  reg [32-1:0] conv2d_25_stream_act_local_5;
  reg [32-1:0] conv2d_25_stream_act_local_6;
  reg [32-1:0] conv2d_25_stream_act_local_7;
  reg [32-1:0] conv2d_25_stream_act_local_8;
  reg [32-1:0] conv2d_25_stream_out_local_val;
  reg [32-1:0] conv2d_25_stream_out_local_col;
  wire [32-1:0] conv2d_25_stream_out_local;
  assign conv2d_25_stream_out_local = conv2d_25_stream_out_local_val + conv2d_25_stream_out_local_col;
  reg [32-1:0] conv2d_25_act_page_comp_offset_0;
  reg [32-1:0] conv2d_25_act_page_comp_offset_1;
  reg [32-1:0] conv2d_25_act_page_comp_offset_2;
  reg [32-1:0] conv2d_25_act_page_dma_offset_0;
  reg [32-1:0] conv2d_25_act_page_dma_offset_1;
  reg [32-1:0] conv2d_25_act_page_dma_offset_2;
  reg [32-1:0] conv2d_25_filter_page_comp_offset;
  reg [32-1:0] conv2d_25_filter_page_dma_offset;
  reg conv2d_25_out_page;
  reg [32-1:0] conv2d_25_out_page_comp_offset;
  reg [32-1:0] conv2d_25_out_page_dma_offset;
  reg [32-1:0] conv2d_25_out_laddr_offset;
  reg conv2d_25_skip_read_filter;
  reg conv2d_25_skip_read_act;
  reg conv2d_25_skip_comp;
  reg conv2d_25_skip_write_out;
  wire [32-1:0] mask_addr_shifted_54;
  assign mask_addr_shifted_54 = conv2d_25_arg_objaddr_2 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_55;
  assign mask_addr_masked_55 = mask_addr_shifted_54 << 2;
  reg [32-1:0] _maxi_read_req_fsm;
  localparam _maxi_read_req_fsm_init = 0;
  reg [33-1:0] _maxi_read_cur_global_size;
  reg _maxi_read_cont;
  wire [8-1:0] pack_read_req_op_sel_56;
  wire [32-1:0] pack_read_req_local_addr_57;
  wire [32-1:0] pack_read_req_local_stride_58;
  wire [33-1:0] pack_read_req_local_size_59;
  wire [32-1:0] pack_read_req_local_blocksize_60;
  assign pack_read_req_op_sel_56 = _maxi_read_op_sel;
  assign pack_read_req_local_addr_57 = _maxi_read_local_addr;
  assign pack_read_req_local_stride_58 = _maxi_read_local_stride;
  assign pack_read_req_local_size_59 = _maxi_read_local_size;
  assign pack_read_req_local_blocksize_60 = _maxi_read_local_blocksize;
  wire [137-1:0] pack_read_req_packed_61;
  assign pack_read_req_packed_61 = { pack_read_req_op_sel_56, pack_read_req_local_addr_57, pack_read_req_local_stride_58, pack_read_req_local_size_59, pack_read_req_local_blocksize_60 };
  assign _maxi_read_req_fifo_wdata = ((_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full)? pack_read_req_packed_61 : 'hx;
  assign _maxi_read_req_fifo_enq = ((_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full)? (_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full && !_maxi_read_req_fifo_almost_full : 0;
  localparam _tmp_62 = 1;
  wire [_tmp_62-1:0] _tmp_63;
  assign _tmp_63 = !_maxi_read_req_fifo_almost_full;
  reg [_tmp_62-1:0] __tmp_63_1;
  wire [32-1:0] mask_addr_shifted_64;
  assign mask_addr_shifted_64 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_65;
  assign mask_addr_masked_65 = mask_addr_shifted_64 << 2;
  wire [32-1:0] mask_addr_shifted_66;
  assign mask_addr_shifted_66 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_67;
  assign mask_addr_masked_67 = mask_addr_shifted_66 << 2;
  wire [32-1:0] mask_addr_shifted_68;
  assign mask_addr_shifted_68 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_69;
  assign mask_addr_masked_69 = mask_addr_shifted_68 << 2;
  wire [32-1:0] mask_addr_shifted_70;
  assign mask_addr_shifted_70 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_71;
  assign mask_addr_masked_71 = mask_addr_shifted_70 << 2;
  wire [32-1:0] mask_addr_shifted_72;
  assign mask_addr_shifted_72 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_73;
  assign mask_addr_masked_73 = mask_addr_shifted_72 << 2;
  wire [32-1:0] mask_addr_shifted_74;
  assign mask_addr_shifted_74 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_75;
  assign mask_addr_masked_75 = mask_addr_shifted_74 << 2;
  reg _maxi_raddr_cond_0_1;
  reg [32-1:0] _maxi_read_data_fsm;
  localparam _maxi_read_data_fsm_init = 0;
  reg [32-1:0] write_burst_fsm_0;
  localparam write_burst_fsm_0_init = 0;
  reg [12-1:0] write_burst_addr_76;
  reg [12-1:0] write_burst_stride_77;
  reg [33-1:0] write_burst_length_78;
  reg write_burst_done_79;
  assign ram_w32_l4096_id0_1_addr = ((write_burst_fsm_0 == 1) && _maxi_rvalid_sb_0)? write_burst_addr_76 : 'hx;
  assign ram_w32_l4096_id0_1_wdata = ((write_burst_fsm_0 == 1) && _maxi_rvalid_sb_0)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l4096_id0_1_wenable = ((write_burst_fsm_0 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w32_l4096_id0_1_enable = ((write_burst_fsm_0 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [32-1:0] mask_addr_shifted_80;
  assign mask_addr_shifted_80 = conv2d_25_arg_objaddr_3 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_81;
  assign mask_addr_masked_81 = mask_addr_shifted_80 << 2;
  reg [32-1:0] write_burst_fsm_1;
  localparam write_burst_fsm_1_init = 0;
  reg [10-1:0] write_burst_addr_82;
  reg [10-1:0] write_burst_stride_83;
  reg [33-1:0] write_burst_length_84;
  reg write_burst_done_85;
  assign ram_w32_l1024_id0_1_addr = ((write_burst_fsm_1 == 1) && _maxi_rvalid_sb_0)? write_burst_addr_82 : 'hx;
  assign ram_w32_l1024_id0_1_wdata = ((write_burst_fsm_1 == 1) && _maxi_rvalid_sb_0)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l1024_id0_1_wenable = ((write_burst_fsm_1 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w32_l1024_id0_1_enable = ((write_burst_fsm_1 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [32-1:0] mask_addr_shifted_86;
  assign mask_addr_shifted_86 = conv2d_25_arg_objaddr_1 + conv2d_25_filter_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_87;
  assign mask_addr_masked_87 = mask_addr_shifted_86 << 2;
  wire write_burst_block_ram_wvalid_88;
  wire write_burst_block_ram_wquit_89;
  reg [32-1:0] write_burst_fsm_2;
  localparam write_burst_fsm_2_init = 0;
  reg [10-1:0] write_burst_addr_90;
  reg [10-1:0] write_burst_stride_91;
  reg [33-1:0] write_burst_length_92;
  reg write_burst_done_93;
  assign ram_w32_l1024_id2_1_addr = ((write_burst_fsm_2 == 1) && write_burst_block_ram_wvalid_88)? write_burst_addr_90 : 'hx;
  assign ram_w32_l1024_id2_1_wdata = ((write_burst_fsm_2 == 1) && write_burst_block_ram_wvalid_88)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l1024_id2_1_wenable = ((write_burst_fsm_2 == 1) && write_burst_block_ram_wvalid_88)? 1'd1 : 0;
  assign ram_w32_l1024_id2_1_enable = ((write_burst_fsm_2 == 1) && write_burst_block_ram_wvalid_88)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_94;
  wire write_burst_block_ram_wquit_95;
  reg [32-1:0] write_burst_fsm_3;
  localparam write_burst_fsm_3_init = 0;
  reg [10-1:0] write_burst_addr_96;
  reg [10-1:0] write_burst_stride_97;
  reg [33-1:0] write_burst_length_98;
  reg write_burst_done_99;
  assign ram_w32_l1024_id3_1_addr = ((write_burst_fsm_3 == 1) && write_burst_block_ram_wvalid_94)? write_burst_addr_96 : 'hx;
  assign ram_w32_l1024_id3_1_wdata = ((write_burst_fsm_3 == 1) && write_burst_block_ram_wvalid_94)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l1024_id3_1_wenable = ((write_burst_fsm_3 == 1) && write_burst_block_ram_wvalid_94)? 1'd1 : 0;
  assign ram_w32_l1024_id3_1_enable = ((write_burst_fsm_3 == 1) && write_burst_block_ram_wvalid_94)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_100;
  wire write_burst_block_ram_wquit_101;
  reg [32-1:0] write_burst_fsm_4;
  localparam write_burst_fsm_4_init = 0;
  reg [10-1:0] write_burst_addr_102;
  reg [10-1:0] write_burst_stride_103;
  reg [33-1:0] write_burst_length_104;
  reg write_burst_done_105;
  assign ram_w32_l1024_id4_1_addr = ((write_burst_fsm_4 == 1) && write_burst_block_ram_wvalid_100)? write_burst_addr_102 : 'hx;
  assign ram_w32_l1024_id4_1_wdata = ((write_burst_fsm_4 == 1) && write_burst_block_ram_wvalid_100)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l1024_id4_1_wenable = ((write_burst_fsm_4 == 1) && write_burst_block_ram_wvalid_100)? 1'd1 : 0;
  assign ram_w32_l1024_id4_1_enable = ((write_burst_fsm_4 == 1) && write_burst_block_ram_wvalid_100)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_106;
  wire write_burst_block_ram_wquit_107;
  reg [32-1:0] write_burst_fsm_5;
  localparam write_burst_fsm_5_init = 0;
  reg [10-1:0] write_burst_addr_108;
  reg [10-1:0] write_burst_stride_109;
  reg [33-1:0] write_burst_length_110;
  reg write_burst_done_111;
  assign ram_w32_l1024_id5_1_addr = ((write_burst_fsm_5 == 1) && write_burst_block_ram_wvalid_106)? write_burst_addr_108 : 'hx;
  assign ram_w32_l1024_id5_1_wdata = ((write_burst_fsm_5 == 1) && write_burst_block_ram_wvalid_106)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l1024_id5_1_wenable = ((write_burst_fsm_5 == 1) && write_burst_block_ram_wvalid_106)? 1'd1 : 0;
  assign ram_w32_l1024_id5_1_enable = ((write_burst_fsm_5 == 1) && write_burst_block_ram_wvalid_106)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_112;
  wire write_burst_block_ram_wquit_113;
  reg [32-1:0] write_burst_fsm_6;
  localparam write_burst_fsm_6_init = 0;
  reg [10-1:0] write_burst_addr_114;
  reg [10-1:0] write_burst_stride_115;
  reg [33-1:0] write_burst_length_116;
  reg write_burst_done_117;
  assign ram_w32_l1024_id6_1_addr = ((write_burst_fsm_6 == 1) && write_burst_block_ram_wvalid_112)? write_burst_addr_114 : 'hx;
  assign ram_w32_l1024_id6_1_wdata = ((write_burst_fsm_6 == 1) && write_burst_block_ram_wvalid_112)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l1024_id6_1_wenable = ((write_burst_fsm_6 == 1) && write_burst_block_ram_wvalid_112)? 1'd1 : 0;
  assign ram_w32_l1024_id6_1_enable = ((write_burst_fsm_6 == 1) && write_burst_block_ram_wvalid_112)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_118;
  wire write_burst_block_ram_wquit_119;
  reg [32-1:0] write_burst_fsm_7;
  localparam write_burst_fsm_7_init = 0;
  reg [10-1:0] write_burst_addr_120;
  reg [10-1:0] write_burst_stride_121;
  reg [33-1:0] write_burst_length_122;
  reg write_burst_done_123;
  assign ram_w32_l1024_id7_1_addr = ((write_burst_fsm_7 == 1) && write_burst_block_ram_wvalid_118)? write_burst_addr_120 : 'hx;
  assign ram_w32_l1024_id7_1_wdata = ((write_burst_fsm_7 == 1) && write_burst_block_ram_wvalid_118)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l1024_id7_1_wenable = ((write_burst_fsm_7 == 1) && write_burst_block_ram_wvalid_118)? 1'd1 : 0;
  assign ram_w32_l1024_id7_1_enable = ((write_burst_fsm_7 == 1) && write_burst_block_ram_wvalid_118)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_124;
  wire write_burst_block_ram_wquit_125;
  reg [32-1:0] write_burst_fsm_8;
  localparam write_burst_fsm_8_init = 0;
  reg [10-1:0] write_burst_addr_126;
  reg [10-1:0] write_burst_stride_127;
  reg [33-1:0] write_burst_length_128;
  reg write_burst_done_129;
  assign ram_w32_l1024_id8_1_addr = ((write_burst_fsm_8 == 1) && write_burst_block_ram_wvalid_124)? write_burst_addr_126 : 'hx;
  assign ram_w32_l1024_id8_1_wdata = ((write_burst_fsm_8 == 1) && write_burst_block_ram_wvalid_124)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l1024_id8_1_wenable = ((write_burst_fsm_8 == 1) && write_burst_block_ram_wvalid_124)? 1'd1 : 0;
  assign ram_w32_l1024_id8_1_enable = ((write_burst_fsm_8 == 1) && write_burst_block_ram_wvalid_124)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_130;
  wire write_burst_block_ram_wquit_131;
  reg [32-1:0] write_burst_fsm_9;
  localparam write_burst_fsm_9_init = 0;
  reg [10-1:0] write_burst_addr_132;
  reg [10-1:0] write_burst_stride_133;
  reg [33-1:0] write_burst_length_134;
  reg write_burst_done_135;
  assign ram_w32_l1024_id9_1_addr = ((write_burst_fsm_9 == 1) && write_burst_block_ram_wvalid_130)? write_burst_addr_132 : 'hx;
  assign ram_w32_l1024_id9_1_wdata = ((write_burst_fsm_9 == 1) && write_burst_block_ram_wvalid_130)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l1024_id9_1_wenable = ((write_burst_fsm_9 == 1) && write_burst_block_ram_wvalid_130)? 1'd1 : 0;
  assign ram_w32_l1024_id9_1_enable = ((write_burst_fsm_9 == 1) && write_burst_block_ram_wvalid_130)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_136;
  wire write_burst_block_ram_wquit_137;
  reg [32-1:0] write_burst_fsm_10;
  localparam write_burst_fsm_10_init = 0;
  reg [10-1:0] write_burst_addr_138;
  reg [10-1:0] write_burst_stride_139;
  reg [33-1:0] write_burst_length_140;
  reg write_burst_done_141;
  assign ram_w32_l1024_id10_1_addr = ((write_burst_fsm_10 == 1) && write_burst_block_ram_wvalid_136)? write_burst_addr_138 : 'hx;
  assign ram_w32_l1024_id10_1_wdata = ((write_burst_fsm_10 == 1) && write_burst_block_ram_wvalid_136)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l1024_id10_1_wenable = ((write_burst_fsm_10 == 1) && write_burst_block_ram_wvalid_136)? 1'd1 : 0;
  assign ram_w32_l1024_id10_1_enable = ((write_burst_fsm_10 == 1) && write_burst_block_ram_wvalid_136)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_11;
  localparam write_burst_block_fsm_11_init = 0;
  reg [33-1:0] write_burst_block_length_142;
  reg [32-1:0] write_burst_block_blocksize_143;
  reg write_burst_block_done_144;
  reg [32-1:0] write_burst_block_count_145;
  assign write_burst_block_ram_wvalid_88 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 1);
  assign write_burst_block_ram_wquit_89 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1);
  assign write_burst_block_ram_wvalid_94 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 2);
  assign write_burst_block_ram_wquit_95 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1);
  assign write_burst_block_ram_wvalid_100 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 3);
  assign write_burst_block_ram_wquit_101 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1);
  assign write_burst_block_ram_wvalid_106 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 4);
  assign write_burst_block_ram_wquit_107 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1);
  assign write_burst_block_ram_wvalid_112 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 5);
  assign write_burst_block_ram_wquit_113 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1);
  assign write_burst_block_ram_wvalid_118 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 6);
  assign write_burst_block_ram_wquit_119 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1);
  assign write_burst_block_ram_wvalid_124 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 7);
  assign write_burst_block_ram_wquit_125 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1);
  assign write_burst_block_ram_wvalid_130 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 8);
  assign write_burst_block_ram_wquit_131 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1);
  assign write_burst_block_ram_wvalid_136 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 9);
  assign write_burst_block_ram_wquit_137 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1);
  wire [32-1:0] conv2d_25_mux_act_gaddr_0;
  assign conv2d_25_mux_act_gaddr_0 = (conv2d_25_row_select == 0)? conv2d_25_arg_objaddr_0 + (conv2d_25_act_base_offset + cparam_conv2d_25_act_offset_values_0) : 
                                     (conv2d_25_row_select == 1)? conv2d_25_arg_objaddr_0 + (conv2d_25_act_base_offset + cparam_conv2d_25_act_offset_values_2) : 
                                     (conv2d_25_row_select == 2)? conv2d_25_arg_objaddr_0 + (conv2d_25_act_base_offset + cparam_conv2d_25_act_offset_values_1) : 1'd0;
  wire [32-1:0] conv2d_25_mux_act_gaddr_1;
  assign conv2d_25_mux_act_gaddr_1 = (conv2d_25_row_select == 0)? conv2d_25_arg_objaddr_0 + (conv2d_25_act_base_offset + cparam_conv2d_25_act_offset_values_1) : 
                                     (conv2d_25_row_select == 1)? conv2d_25_arg_objaddr_0 + (conv2d_25_act_base_offset + cparam_conv2d_25_act_offset_values_0) : 
                                     (conv2d_25_row_select == 2)? conv2d_25_arg_objaddr_0 + (conv2d_25_act_base_offset + cparam_conv2d_25_act_offset_values_2) : 1'd0;
  wire [32-1:0] conv2d_25_mux_act_gaddr_2;
  assign conv2d_25_mux_act_gaddr_2 = (conv2d_25_row_select == 0)? conv2d_25_arg_objaddr_0 + (conv2d_25_act_base_offset + cparam_conv2d_25_act_offset_values_2) : 
                                     (conv2d_25_row_select == 1)? conv2d_25_arg_objaddr_0 + (conv2d_25_act_base_offset + cparam_conv2d_25_act_offset_values_1) : 
                                     (conv2d_25_row_select == 2)? conv2d_25_arg_objaddr_0 + (conv2d_25_act_base_offset + cparam_conv2d_25_act_offset_values_0) : 1'd0;
  wire conv2d_25_dma_pad_mask_0;
  assign conv2d_25_dma_pad_mask_0 = (conv2d_25_row_count + 0 < cparam_conv2d_25_pad_row_top) || (conv2d_25_row_count + 0 >= cparam_conv2d_25_act_num_row + cparam_conv2d_25_pad_row_top);
  wire conv2d_25_dma_pad_mask_1;
  assign conv2d_25_dma_pad_mask_1 = (conv2d_25_row_count + 1 < cparam_conv2d_25_pad_row_top) || (conv2d_25_row_count + 1 >= cparam_conv2d_25_act_num_row + cparam_conv2d_25_pad_row_top);
  wire conv2d_25_dma_pad_mask_2;
  assign conv2d_25_dma_pad_mask_2 = (conv2d_25_row_count + 2 < cparam_conv2d_25_pad_row_top) || (conv2d_25_row_count + 2 >= cparam_conv2d_25_act_num_row + cparam_conv2d_25_pad_row_top);
  wire conv2d_25_mux_dma_pad_mask_0;
  assign conv2d_25_mux_dma_pad_mask_0 = (conv2d_25_row_select == 0)? conv2d_25_dma_pad_mask_0 : 
                                        (conv2d_25_row_select == 1)? conv2d_25_dma_pad_mask_2 : 
                                        (conv2d_25_row_select == 2)? conv2d_25_dma_pad_mask_1 : 1'd0;
  wire conv2d_25_mux_dma_pad_mask_1;
  assign conv2d_25_mux_dma_pad_mask_1 = (conv2d_25_row_select == 0)? conv2d_25_dma_pad_mask_1 : 
                                        (conv2d_25_row_select == 1)? conv2d_25_dma_pad_mask_0 : 
                                        (conv2d_25_row_select == 2)? conv2d_25_dma_pad_mask_2 : 1'd0;
  wire conv2d_25_mux_dma_pad_mask_2;
  assign conv2d_25_mux_dma_pad_mask_2 = (conv2d_25_row_select == 0)? conv2d_25_dma_pad_mask_2 : 
                                        (conv2d_25_row_select == 1)? conv2d_25_dma_pad_mask_1 : 
                                        (conv2d_25_row_select == 2)? conv2d_25_dma_pad_mask_0 : 1'd0;
  wire conv2d_25_mux_dma_flag_0;
  assign conv2d_25_mux_dma_flag_0 = (conv2d_25_prev_row_select == 0)? conv2d_25_dma_flag_0 : 
                                    (conv2d_25_prev_row_select == 1)? conv2d_25_dma_flag_2 : 
                                    (conv2d_25_prev_row_select == 2)? conv2d_25_dma_flag_1 : 1'd0;
  wire conv2d_25_mux_dma_flag_1;
  assign conv2d_25_mux_dma_flag_1 = (conv2d_25_prev_row_select == 0)? conv2d_25_dma_flag_1 : 
                                    (conv2d_25_prev_row_select == 1)? conv2d_25_dma_flag_0 : 
                                    (conv2d_25_prev_row_select == 2)? conv2d_25_dma_flag_2 : 1'd0;
  wire conv2d_25_mux_dma_flag_2;
  assign conv2d_25_mux_dma_flag_2 = (conv2d_25_prev_row_select == 0)? conv2d_25_dma_flag_2 : 
                                    (conv2d_25_prev_row_select == 1)? conv2d_25_dma_flag_1 : 
                                    (conv2d_25_prev_row_select == 2)? conv2d_25_dma_flag_0 : 1'd0;
  wire [32-1:0] mask_addr_shifted_146;
  assign mask_addr_shifted_146 = conv2d_25_mux_act_gaddr_0 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_147;
  assign mask_addr_masked_147 = mask_addr_shifted_146 << 2;
  wire write_burst_block_ram_wvalid_148;
  wire write_burst_block_ram_wquit_149;
  reg [32-1:0] write_burst_fsm_12;
  localparam write_burst_fsm_12_init = 0;
  reg [12-1:0] write_burst_addr_150;
  reg [12-1:0] write_burst_stride_151;
  reg [33-1:0] write_burst_length_152;
  reg write_burst_done_153;
  assign ram_w32_l4096_id1_1_addr = ((write_burst_fsm_12 == 1) && write_burst_block_ram_wvalid_148)? write_burst_addr_150 : 'hx;
  assign ram_w32_l4096_id1_1_wdata = ((write_burst_fsm_12 == 1) && write_burst_block_ram_wvalid_148)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l4096_id1_1_wenable = ((write_burst_fsm_12 == 1) && write_burst_block_ram_wvalid_148)? 1'd1 : 0;
  assign ram_w32_l4096_id1_1_enable = ((write_burst_fsm_12 == 1) && write_burst_block_ram_wvalid_148)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_154;
  wire write_burst_block_ram_wquit_155;
  reg [32-1:0] write_burst_fsm_13;
  localparam write_burst_fsm_13_init = 0;
  reg [12-1:0] write_burst_addr_156;
  reg [12-1:0] write_burst_stride_157;
  reg [33-1:0] write_burst_length_158;
  reg write_burst_done_159;
  assign ram_w32_l4096_id2_1_addr = ((write_burst_fsm_13 == 1) && write_burst_block_ram_wvalid_154)? write_burst_addr_156 : 'hx;
  assign ram_w32_l4096_id2_1_wdata = ((write_burst_fsm_13 == 1) && write_burst_block_ram_wvalid_154)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l4096_id2_1_wenable = ((write_burst_fsm_13 == 1) && write_burst_block_ram_wvalid_154)? 1'd1 : 0;
  assign ram_w32_l4096_id2_1_enable = ((write_burst_fsm_13 == 1) && write_burst_block_ram_wvalid_154)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_160;
  wire write_burst_block_ram_wquit_161;
  reg [32-1:0] write_burst_fsm_14;
  localparam write_burst_fsm_14_init = 0;
  reg [12-1:0] write_burst_addr_162;
  reg [12-1:0] write_burst_stride_163;
  reg [33-1:0] write_burst_length_164;
  reg write_burst_done_165;
  assign ram_w32_l4096_id3_1_addr = ((write_burst_fsm_14 == 1) && write_burst_block_ram_wvalid_160)? write_burst_addr_162 : 'hx;
  assign ram_w32_l4096_id3_1_wdata = ((write_burst_fsm_14 == 1) && write_burst_block_ram_wvalid_160)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l4096_id3_1_wenable = ((write_burst_fsm_14 == 1) && write_burst_block_ram_wvalid_160)? 1'd1 : 0;
  assign ram_w32_l4096_id3_1_enable = ((write_burst_fsm_14 == 1) && write_burst_block_ram_wvalid_160)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_15;
  localparam write_burst_block_fsm_15_init = 0;
  reg [33-1:0] write_burst_block_length_166;
  reg [32-1:0] write_burst_block_blocksize_167;
  reg write_burst_block_done_168;
  reg [32-1:0] write_burst_block_count_169;
  assign write_burst_block_ram_wvalid_148 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_15 == 1);
  assign write_burst_block_ram_wquit_149 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_166 <= 1);
  assign write_burst_block_ram_wvalid_154 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_15 == 2);
  assign write_burst_block_ram_wquit_155 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_166 <= 1);
  assign write_burst_block_ram_wvalid_160 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_15 == 3);
  assign write_burst_block_ram_wquit_161 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_166 <= 1);
  wire [32-1:0] mask_addr_shifted_170;
  assign mask_addr_shifted_170 = conv2d_25_mux_act_gaddr_1 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_171;
  assign mask_addr_masked_171 = mask_addr_shifted_170 << 2;
  wire write_burst_block_ram_wvalid_172;
  wire write_burst_block_ram_wquit_173;
  reg [32-1:0] write_burst_fsm_16;
  localparam write_burst_fsm_16_init = 0;
  reg [12-1:0] write_burst_addr_174;
  reg [12-1:0] write_burst_stride_175;
  reg [33-1:0] write_burst_length_176;
  reg write_burst_done_177;
  assign ram_w32_l4096_id4_1_addr = ((write_burst_fsm_16 == 1) && write_burst_block_ram_wvalid_172)? write_burst_addr_174 : 'hx;
  assign ram_w32_l4096_id4_1_wdata = ((write_burst_fsm_16 == 1) && write_burst_block_ram_wvalid_172)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l4096_id4_1_wenable = ((write_burst_fsm_16 == 1) && write_burst_block_ram_wvalid_172)? 1'd1 : 0;
  assign ram_w32_l4096_id4_1_enable = ((write_burst_fsm_16 == 1) && write_burst_block_ram_wvalid_172)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_178;
  wire write_burst_block_ram_wquit_179;
  reg [32-1:0] write_burst_fsm_17;
  localparam write_burst_fsm_17_init = 0;
  reg [12-1:0] write_burst_addr_180;
  reg [12-1:0] write_burst_stride_181;
  reg [33-1:0] write_burst_length_182;
  reg write_burst_done_183;
  assign ram_w32_l4096_id5_1_addr = ((write_burst_fsm_17 == 1) && write_burst_block_ram_wvalid_178)? write_burst_addr_180 : 'hx;
  assign ram_w32_l4096_id5_1_wdata = ((write_burst_fsm_17 == 1) && write_burst_block_ram_wvalid_178)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l4096_id5_1_wenable = ((write_burst_fsm_17 == 1) && write_burst_block_ram_wvalid_178)? 1'd1 : 0;
  assign ram_w32_l4096_id5_1_enable = ((write_burst_fsm_17 == 1) && write_burst_block_ram_wvalid_178)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_184;
  wire write_burst_block_ram_wquit_185;
  reg [32-1:0] write_burst_fsm_18;
  localparam write_burst_fsm_18_init = 0;
  reg [12-1:0] write_burst_addr_186;
  reg [12-1:0] write_burst_stride_187;
  reg [33-1:0] write_burst_length_188;
  reg write_burst_done_189;
  assign ram_w32_l4096_id6_1_addr = ((write_burst_fsm_18 == 1) && write_burst_block_ram_wvalid_184)? write_burst_addr_186 : 'hx;
  assign ram_w32_l4096_id6_1_wdata = ((write_burst_fsm_18 == 1) && write_burst_block_ram_wvalid_184)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l4096_id6_1_wenable = ((write_burst_fsm_18 == 1) && write_burst_block_ram_wvalid_184)? 1'd1 : 0;
  assign ram_w32_l4096_id6_1_enable = ((write_burst_fsm_18 == 1) && write_burst_block_ram_wvalid_184)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_19;
  localparam write_burst_block_fsm_19_init = 0;
  reg [33-1:0] write_burst_block_length_190;
  reg [32-1:0] write_burst_block_blocksize_191;
  reg write_burst_block_done_192;
  reg [32-1:0] write_burst_block_count_193;
  assign write_burst_block_ram_wvalid_172 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_19 == 1);
  assign write_burst_block_ram_wquit_173 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_190 <= 1);
  assign write_burst_block_ram_wvalid_178 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_19 == 2);
  assign write_burst_block_ram_wquit_179 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_190 <= 1);
  assign write_burst_block_ram_wvalid_184 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_19 == 3);
  assign write_burst_block_ram_wquit_185 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_190 <= 1);
  wire [32-1:0] mask_addr_shifted_194;
  assign mask_addr_shifted_194 = conv2d_25_mux_act_gaddr_2 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_195;
  assign mask_addr_masked_195 = mask_addr_shifted_194 << 2;
  wire write_burst_block_ram_wvalid_196;
  wire write_burst_block_ram_wquit_197;
  reg [32-1:0] write_burst_fsm_20;
  localparam write_burst_fsm_20_init = 0;
  reg [12-1:0] write_burst_addr_198;
  reg [12-1:0] write_burst_stride_199;
  reg [33-1:0] write_burst_length_200;
  reg write_burst_done_201;
  assign ram_w32_l4096_id7_1_addr = ((write_burst_fsm_20 == 1) && write_burst_block_ram_wvalid_196)? write_burst_addr_198 : 'hx;
  assign ram_w32_l4096_id7_1_wdata = ((write_burst_fsm_20 == 1) && write_burst_block_ram_wvalid_196)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l4096_id7_1_wenable = ((write_burst_fsm_20 == 1) && write_burst_block_ram_wvalid_196)? 1'd1 : 0;
  assign ram_w32_l4096_id7_1_enable = ((write_burst_fsm_20 == 1) && write_burst_block_ram_wvalid_196)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_202;
  wire write_burst_block_ram_wquit_203;
  reg [32-1:0] write_burst_fsm_21;
  localparam write_burst_fsm_21_init = 0;
  reg [12-1:0] write_burst_addr_204;
  reg [12-1:0] write_burst_stride_205;
  reg [33-1:0] write_burst_length_206;
  reg write_burst_done_207;
  assign ram_w32_l4096_id8_1_addr = ((write_burst_fsm_21 == 1) && write_burst_block_ram_wvalid_202)? write_burst_addr_204 : 'hx;
  assign ram_w32_l4096_id8_1_wdata = ((write_burst_fsm_21 == 1) && write_burst_block_ram_wvalid_202)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l4096_id8_1_wenable = ((write_burst_fsm_21 == 1) && write_burst_block_ram_wvalid_202)? 1'd1 : 0;
  assign ram_w32_l4096_id8_1_enable = ((write_burst_fsm_21 == 1) && write_burst_block_ram_wvalid_202)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_208;
  wire write_burst_block_ram_wquit_209;
  reg [32-1:0] write_burst_fsm_22;
  localparam write_burst_fsm_22_init = 0;
  reg [13-1:0] write_burst_addr_210;
  reg [13-1:0] write_burst_stride_211;
  reg [33-1:0] write_burst_length_212;
  reg write_burst_done_213;
  reg [32-1:0] write_burst_block_fsm_23;
  localparam write_burst_block_fsm_23_init = 0;
  reg [33-1:0] write_burst_block_length_214;
  reg [32-1:0] write_burst_block_blocksize_215;
  reg write_burst_block_done_216;
  reg [32-1:0] write_burst_block_count_217;
  assign write_burst_block_ram_wvalid_196 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_23 == 1);
  assign write_burst_block_ram_wquit_197 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_214 <= 1);
  assign write_burst_block_ram_wvalid_202 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_23 == 2);
  assign write_burst_block_ram_wquit_203 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_214 <= 1);
  assign write_burst_block_ram_wvalid_208 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_23 == 3);
  assign write_burst_block_ram_wquit_209 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_214 <= 1);
  reg [32-1:0] conv2d_25_comp_fsm;
  localparam conv2d_25_comp_fsm_init = 0;
  reg [32-1:0] conv2d_25_filter_page_comp_offset_buf;
  reg [32-1:0] conv2d_25_act_page_comp_offset_buf_0;
  reg [32-1:0] conv2d_25_act_page_comp_offset_buf_1;
  reg [32-1:0] conv2d_25_act_page_comp_offset_buf_2;
  reg [32-1:0] conv2d_25_out_page_comp_offset_buf;
  reg [32-1:0] conv2d_25_row_count_buf;
  reg [2-1:0] conv2d_25_row_select_buf;
  reg [32-1:0] conv2d_25_och_count_buf;
  wire conv2d_25_stream_pad_mask_0_0;
  assign conv2d_25_stream_pad_mask_0_0 = (conv2d_25_col_count + 0 < cparam_conv2d_25_pad_col_left) || (conv2d_25_col_count + 0 >= cparam_conv2d_25_act_num_col + cparam_conv2d_25_pad_col_left) || (conv2d_25_row_count_buf + 0 < cparam_conv2d_25_pad_row_top) || (conv2d_25_row_count_buf + 0 >= cparam_conv2d_25_act_num_row + cparam_conv2d_25_pad_row_top);
  wire conv2d_25_stream_pad_mask_0_1;
  assign conv2d_25_stream_pad_mask_0_1 = (conv2d_25_col_count + 1 < cparam_conv2d_25_pad_col_left) || (conv2d_25_col_count + 1 >= cparam_conv2d_25_act_num_col + cparam_conv2d_25_pad_col_left) || (conv2d_25_row_count_buf + 0 < cparam_conv2d_25_pad_row_top) || (conv2d_25_row_count_buf + 0 >= cparam_conv2d_25_act_num_row + cparam_conv2d_25_pad_row_top);
  wire conv2d_25_stream_pad_mask_0_2;
  assign conv2d_25_stream_pad_mask_0_2 = (conv2d_25_col_count + 2 < cparam_conv2d_25_pad_col_left) || (conv2d_25_col_count + 2 >= cparam_conv2d_25_act_num_col + cparam_conv2d_25_pad_col_left) || (conv2d_25_row_count_buf + 0 < cparam_conv2d_25_pad_row_top) || (conv2d_25_row_count_buf + 0 >= cparam_conv2d_25_act_num_row + cparam_conv2d_25_pad_row_top);
  wire conv2d_25_stream_pad_mask_1_0;
  assign conv2d_25_stream_pad_mask_1_0 = (conv2d_25_col_count + 0 < cparam_conv2d_25_pad_col_left) || (conv2d_25_col_count + 0 >= cparam_conv2d_25_act_num_col + cparam_conv2d_25_pad_col_left) || (conv2d_25_row_count_buf + 1 < cparam_conv2d_25_pad_row_top) || (conv2d_25_row_count_buf + 1 >= cparam_conv2d_25_act_num_row + cparam_conv2d_25_pad_row_top);
  wire conv2d_25_stream_pad_mask_1_1;
  assign conv2d_25_stream_pad_mask_1_1 = (conv2d_25_col_count + 1 < cparam_conv2d_25_pad_col_left) || (conv2d_25_col_count + 1 >= cparam_conv2d_25_act_num_col + cparam_conv2d_25_pad_col_left) || (conv2d_25_row_count_buf + 1 < cparam_conv2d_25_pad_row_top) || (conv2d_25_row_count_buf + 1 >= cparam_conv2d_25_act_num_row + cparam_conv2d_25_pad_row_top);
  wire conv2d_25_stream_pad_mask_1_2;
  assign conv2d_25_stream_pad_mask_1_2 = (conv2d_25_col_count + 2 < cparam_conv2d_25_pad_col_left) || (conv2d_25_col_count + 2 >= cparam_conv2d_25_act_num_col + cparam_conv2d_25_pad_col_left) || (conv2d_25_row_count_buf + 1 < cparam_conv2d_25_pad_row_top) || (conv2d_25_row_count_buf + 1 >= cparam_conv2d_25_act_num_row + cparam_conv2d_25_pad_row_top);
  wire conv2d_25_stream_pad_mask_2_0;
  assign conv2d_25_stream_pad_mask_2_0 = (conv2d_25_col_count + 0 < cparam_conv2d_25_pad_col_left) || (conv2d_25_col_count + 0 >= cparam_conv2d_25_act_num_col + cparam_conv2d_25_pad_col_left) || (conv2d_25_row_count_buf + 2 < cparam_conv2d_25_pad_row_top) || (conv2d_25_row_count_buf + 2 >= cparam_conv2d_25_act_num_row + cparam_conv2d_25_pad_row_top);
  wire conv2d_25_stream_pad_mask_2_1;
  assign conv2d_25_stream_pad_mask_2_1 = (conv2d_25_col_count + 1 < cparam_conv2d_25_pad_col_left) || (conv2d_25_col_count + 1 >= cparam_conv2d_25_act_num_col + cparam_conv2d_25_pad_col_left) || (conv2d_25_row_count_buf + 2 < cparam_conv2d_25_pad_row_top) || (conv2d_25_row_count_buf + 2 >= cparam_conv2d_25_act_num_row + cparam_conv2d_25_pad_row_top);
  wire conv2d_25_stream_pad_mask_2_2;
  assign conv2d_25_stream_pad_mask_2_2 = (conv2d_25_col_count + 2 < cparam_conv2d_25_pad_col_left) || (conv2d_25_col_count + 2 >= cparam_conv2d_25_act_num_col + cparam_conv2d_25_pad_col_left) || (conv2d_25_row_count_buf + 2 < cparam_conv2d_25_pad_row_top) || (conv2d_25_row_count_buf + 2 >= cparam_conv2d_25_act_num_row + cparam_conv2d_25_pad_row_top);
  reg [9-1:0] conv2d_25_stream_pad_masks;
  wire [10-1:0] stream_conv2d_25_parameter_0_data;
  wire [2-1:0] stream_conv2d_25_parameter_1_data;
  wire [2-1:0] stream_conv2d_25_parameter_2_data;
  wire [9-1:0] stream_conv2d_25_parameter_3_data;
  wire [1-1:0] stream_conv2d_25_parameter_4_data;
  wire [1-1:0] stream_conv2d_25__reduce_reset_data;
  wire [1-1:0] stream_conv2d_25_parameter_6_data;
  wire [32-1:0] stream_conv2d_25_source_7_data;
  wire [1-1:0] stream_conv2d_25_parameter_8_data;
  wire [32-1:0] stream_conv2d_25_source_9_data;
  wire [1-1:0] stream_conv2d_25_parameter_10_data;
  wire [32-1:0] stream_conv2d_25_source_11_data;
  wire [1-1:0] stream_conv2d_25_parameter_12_data;
  wire [32-1:0] stream_conv2d_25_source_13_data;
  wire [1-1:0] stream_conv2d_25_parameter_14_data;
  wire [32-1:0] stream_conv2d_25_source_15_data;
  wire [1-1:0] stream_conv2d_25_parameter_16_data;
  wire [1-1:0] stream_conv2d_25_parameter_17_data;
  wire [5-1:0] stream_conv2d_25_parameter_18_data;
  wire [1-1:0] stream_conv2d_25_parameter_19_data;
  wire [32-1:0] stream_conv2d_25_source_20_data;
  wire [32-1:0] stream_conv2d_25_source_21_data;
  wire [32-1:0] stream_conv2d_25_source_22_data;
  wire [32-1:0] stream_conv2d_25_source_23_data;
  wire [32-1:0] stream_conv2d_25_source_24_data;
  wire [32-1:0] stream_conv2d_25_source_25_data;
  wire [32-1:0] stream_conv2d_25_source_26_data;
  wire [32-1:0] stream_conv2d_25_source_27_data;
  wire [32-1:0] stream_conv2d_25_source_28_data;
  wire [32-1:0] stream_conv2d_25_source_29_data;
  wire [32-1:0] stream_conv2d_25_source_30_data;
  wire [32-1:0] stream_conv2d_25_source_31_data;
  wire [32-1:0] stream_conv2d_25_source_32_data;
  wire [32-1:0] stream_conv2d_25_source_33_data;
  wire [32-1:0] stream_conv2d_25_source_34_data;
  wire [32-1:0] stream_conv2d_25_source_35_data;
  wire [32-1:0] stream_conv2d_25_source_36_data;
  wire [32-1:0] stream_conv2d_25_source_37_data;
  reg __stream_conv2d_25_stream_ivalid_1;
  reg __stream_conv2d_25_stream_ivalid_2;
  reg __stream_conv2d_25_stream_ivalid_3;
  reg __stream_conv2d_25_stream_ivalid_4;
  reg __stream_conv2d_25_stream_ivalid_5;
  reg __stream_conv2d_25_stream_ivalid_6;
  reg __stream_conv2d_25_stream_ivalid_7;
  reg __stream_conv2d_25_stream_ivalid_8;
  reg __stream_conv2d_25_stream_ivalid_9;
  reg __stream_conv2d_25_stream_ivalid_10;
  reg __stream_conv2d_25_stream_ivalid_11;
  reg __stream_conv2d_25_stream_ivalid_12;
  reg __stream_conv2d_25_stream_ivalid_13;
  reg __stream_conv2d_25_stream_ivalid_14;
  reg __stream_conv2d_25_stream_ivalid_15;
  reg __stream_conv2d_25_stream_ivalid_16;
  reg __stream_conv2d_25_stream_ivalid_17;
  reg __stream_conv2d_25_stream_ivalid_18;
  reg __stream_conv2d_25_stream_ivalid_19;
  reg __stream_conv2d_25_stream_ivalid_20;
  reg __stream_conv2d_25_stream_ivalid_21;
  reg __stream_conv2d_25_stream_ivalid_22;
  reg __stream_conv2d_25_stream_ivalid_23;
  reg __stream_conv2d_25_stream_ivalid_24;
  reg __stream_conv2d_25_stream_ivalid_25;
  reg __stream_conv2d_25_stream_ivalid_26;
  reg __stream_conv2d_25_stream_ivalid_27;
  reg __stream_conv2d_25_stream_ivalid_28;
  reg __stream_conv2d_25_stream_ivalid_29;
  reg __stream_conv2d_25_stream_ivalid_30;
  reg __stream_conv2d_25_stream_ivalid_31;
  reg __stream_conv2d_25_stream_ivalid_32;
  reg __stream_conv2d_25_stream_ivalid_33;
  reg __stream_conv2d_25_stream_ivalid_34;
  wire [32-1:0] _slice_data_295;
  assign _slice_data_295 = stream_conv2d_25_source_7_data[6'd31:1'd0];
  wire [32-1:0] _reinterpretcast_src_296;
  assign _reinterpretcast_src_296 = _slice_data_295;
  wire signed [32-1:0] _reinterpretcast_data_296;
  assign _reinterpretcast_data_296 = _reinterpretcast_src_296;
  wire signed [32-1:0] _cond_data_297;
  assign _cond_data_297 = (stream_conv2d_25_parameter_6_data)? _reinterpretcast_data_296 : _reinterpretcast_data_296;
  wire [32-1:0] _slice_data_302;
  assign _slice_data_302 = stream_conv2d_25_source_9_data[6'd31:1'd0];
  wire [32-1:0] _reinterpretcast_src_303;
  assign _reinterpretcast_src_303 = _slice_data_302;
  wire signed [32-1:0] _reinterpretcast_data_303;
  assign _reinterpretcast_data_303 = _reinterpretcast_src_303;
  wire signed [32-1:0] _cond_data_304;
  assign _cond_data_304 = (stream_conv2d_25_parameter_8_data)? _reinterpretcast_data_303 : _reinterpretcast_data_303;
  wire [32-1:0] _slice_data_309;
  assign _slice_data_309 = stream_conv2d_25_source_11_data[6'd31:1'd0];
  wire [32-1:0] _reinterpretcast_src_310;
  assign _reinterpretcast_src_310 = _slice_data_309;
  wire [32-1:0] _reinterpretcast_data_310;
  assign _reinterpretcast_data_310 = _reinterpretcast_src_310;
  wire [32-1:0] _cond_data_311;
  assign _cond_data_311 = (stream_conv2d_25_parameter_10_data)? _reinterpretcast_data_310 : _reinterpretcast_data_310;
  wire [32-1:0] _slice_data_316;
  assign _slice_data_316 = stream_conv2d_25_source_13_data[6'd31:1'd0];
  wire [32-1:0] _reinterpretcast_src_317;
  assign _reinterpretcast_src_317 = _slice_data_316;
  wire [32-1:0] _reinterpretcast_data_317;
  assign _reinterpretcast_data_317 = _reinterpretcast_src_317;
  wire [32-1:0] _cond_data_318;
  assign _cond_data_318 = (stream_conv2d_25_parameter_12_data)? _reinterpretcast_data_317 : _reinterpretcast_data_317;
  wire [32-1:0] _slice_data_323;
  assign _slice_data_323 = stream_conv2d_25_source_15_data[6'd31:1'd0];
  wire [32-1:0] _reinterpretcast_src_324;
  assign _reinterpretcast_src_324 = _slice_data_323;
  wire [32-1:0] _reinterpretcast_data_324;
  assign _reinterpretcast_data_324 = _reinterpretcast_src_324;
  wire [32-1:0] _cond_data_325;
  assign _cond_data_325 = (stream_conv2d_25_parameter_14_data)? _reinterpretcast_data_324 : _reinterpretcast_data_324;
  reg [1-1:0] _eq_data_339;
  reg [1-1:0] _eq_data_343;
  reg [1-1:0] _eq_data_346;
  reg [1-1:0] _eq_data_349;
  reg [1-1:0] _eq_data_353;
  reg [1-1:0] _eq_data_356;
  reg [1-1:0] _eq_data_359;
  reg [1-1:0] _eq_data_363;
  reg [1-1:0] _eq_data_366;
  reg [1-1:0] _eq_data_369;
  reg [1-1:0] _eq_data_373;
  reg [1-1:0] _eq_data_376;
  reg [1-1:0] _eq_data_379;
  reg [1-1:0] _eq_data_383;
  reg [1-1:0] _eq_data_386;
  reg [1-1:0] _eq_data_389;
  reg [1-1:0] _eq_data_393;
  reg [1-1:0] _eq_data_396;
  reg [1-1:0] _eq_data_399;
  reg [1-1:0] _eq_data_403;
  reg [1-1:0] _eq_data_406;
  reg [1-1:0] _eq_data_409;
  reg [1-1:0] _eq_data_413;
  reg [1-1:0] _eq_data_416;
  reg [1-1:0] _eq_data_419;
  reg [1-1:0] _eq_data_423;
  reg [1-1:0] _eq_data_426;
  reg [1-1:0] _eq_data_429;
  reg [1-1:0] _eq_data_433;
  reg [1-1:0] _eq_data_436;
  reg [1-1:0] _eq_data_439;
  reg [1-1:0] _eq_data_443;
  reg [1-1:0] _eq_data_446;
  reg [1-1:0] _eq_data_449;
  reg [1-1:0] _eq_data_453;
  reg [1-1:0] _eq_data_456;
  reg [1-1:0] _eq_data_459;
  reg [1-1:0] _eq_data_463;
  reg [1-1:0] _eq_data_466;
  reg [1-1:0] _eq_data_469;
  reg [1-1:0] _eq_data_473;
  reg [1-1:0] _eq_data_476;
  reg [1-1:0] _eq_data_479;
  reg [1-1:0] _eq_data_483;
  reg [1-1:0] _eq_data_486;
  reg [1-1:0] _eq_data_489;
  reg [1-1:0] _eq_data_493;
  reg [1-1:0] _eq_data_496;
  reg [1-1:0] _eq_data_499;
  reg [1-1:0] _eq_data_503;
  reg [1-1:0] _eq_data_506;
  reg [1-1:0] _eq_data_509;
  reg [1-1:0] _eq_data_513;
  reg [1-1:0] _eq_data_516;
  wire [32-1:0] _reinterpretcast_src_609;
  assign _reinterpretcast_src_609 = stream_conv2d_25_source_29_data;
  wire signed [32-1:0] _reinterpretcast_data_609;
  assign _reinterpretcast_data_609 = _reinterpretcast_src_609;
  wire [32-1:0] _reinterpretcast_src_610;
  assign _reinterpretcast_src_610 = stream_conv2d_25_source_30_data;
  wire signed [32-1:0] _reinterpretcast_data_610;
  assign _reinterpretcast_data_610 = _reinterpretcast_src_610;
  wire [32-1:0] _reinterpretcast_src_611;
  assign _reinterpretcast_src_611 = stream_conv2d_25_source_31_data;
  wire signed [32-1:0] _reinterpretcast_data_611;
  assign _reinterpretcast_data_611 = _reinterpretcast_src_611;
  wire [32-1:0] _reinterpretcast_src_612;
  assign _reinterpretcast_src_612 = stream_conv2d_25_source_32_data;
  wire signed [32-1:0] _reinterpretcast_data_612;
  assign _reinterpretcast_data_612 = _reinterpretcast_src_612;
  wire [32-1:0] _reinterpretcast_src_613;
  assign _reinterpretcast_src_613 = stream_conv2d_25_source_33_data;
  wire signed [32-1:0] _reinterpretcast_data_613;
  assign _reinterpretcast_data_613 = _reinterpretcast_src_613;
  wire [32-1:0] _reinterpretcast_src_614;
  assign _reinterpretcast_src_614 = stream_conv2d_25_source_34_data;
  wire signed [32-1:0] _reinterpretcast_data_614;
  assign _reinterpretcast_data_614 = _reinterpretcast_src_614;
  wire [32-1:0] _reinterpretcast_src_615;
  assign _reinterpretcast_src_615 = stream_conv2d_25_source_35_data;
  wire signed [32-1:0] _reinterpretcast_data_615;
  assign _reinterpretcast_data_615 = _reinterpretcast_src_615;
  wire [32-1:0] _reinterpretcast_src_616;
  assign _reinterpretcast_src_616 = stream_conv2d_25_source_36_data;
  wire signed [32-1:0] _reinterpretcast_data_616;
  assign _reinterpretcast_data_616 = _reinterpretcast_src_616;
  wire [32-1:0] _reinterpretcast_src_617;
  assign _reinterpretcast_src_617 = stream_conv2d_25_source_37_data;
  wire signed [32-1:0] _reinterpretcast_data_617;
  assign _reinterpretcast_data_617 = _reinterpretcast_src_617;
  wire [1-1:0] _pointer_data_618;
  assign _pointer_data_618 = stream_conv2d_25_parameter_3_data[1'sd0];
  wire [1-1:0] _pointer_data_620;
  assign _pointer_data_620 = stream_conv2d_25_parameter_3_data[2'sd1];
  wire [1-1:0] _pointer_data_622;
  assign _pointer_data_622 = stream_conv2d_25_parameter_3_data[3'sd2];
  wire [1-1:0] _pointer_data_624;
  assign _pointer_data_624 = stream_conv2d_25_parameter_3_data[3'sd3];
  wire [1-1:0] _pointer_data_626;
  assign _pointer_data_626 = stream_conv2d_25_parameter_3_data[4'sd4];
  wire [1-1:0] _pointer_data_628;
  assign _pointer_data_628 = stream_conv2d_25_parameter_3_data[4'sd5];
  wire [1-1:0] _pointer_data_630;
  assign _pointer_data_630 = stream_conv2d_25_parameter_3_data[4'sd6];
  wire [1-1:0] _pointer_data_632;
  assign _pointer_data_632 = stream_conv2d_25_parameter_3_data[4'sd7];
  wire [1-1:0] _pointer_data_634;
  assign _pointer_data_634 = stream_conv2d_25_parameter_3_data[5'sd8];
  reg [32-1:0] _plus_data_671;
  reg [32-1:0] _plus_data_690;
  reg [32-1:0] _plus_data_709;
  reg [32-1:0] _plus_data_728;
  reg [32-1:0] _plus_data_747;
  reg [32-1:0] _plus_data_766;
  reg [32-1:0] _plus_data_785;
  reg [32-1:0] _plus_data_804;
  reg [32-1:0] _plus_data_823;
  reg [32-1:0] _plus_data_839;
  reg [32-1:0] _plus_data_858;
  wire [1-1:0] _eq_data_873;
  assign _eq_data_873 = 1'sd0 == 6'sd31;
  reg [32-1:0] __delay_data_946__variable_332;
  reg [32-1:0] __delay_data_947__variable_331;
  reg [32-1:0] __delay_data_948__variable_330;
  reg [32-1:0] __delay_data_949__variable_335;
  reg [32-1:0] __delay_data_950__variable_334;
  reg [32-1:0] __delay_data_951__variable_333;
  reg [32-1:0] __delay_data_952__variable_338;
  reg [32-1:0] __delay_data_953__variable_337;
  reg [32-1:0] __delay_data_954__variable_336;
  reg [1-1:0] __delay_data_955_pointer_618;
  reg signed [32-1:0] __delay_data_956_reinterpretcast_609;
  reg [1-1:0] __delay_data_957_pointer_620;
  reg signed [32-1:0] __delay_data_958_reinterpretcast_610;
  reg [1-1:0] __delay_data_959_pointer_622;
  reg signed [32-1:0] __delay_data_960_reinterpretcast_611;
  reg [1-1:0] __delay_data_961_pointer_624;
  reg signed [32-1:0] __delay_data_962_reinterpretcast_612;
  reg [1-1:0] __delay_data_963_pointer_626;
  reg signed [32-1:0] __delay_data_964_reinterpretcast_613;
  reg [1-1:0] __delay_data_965_pointer_628;
  reg signed [32-1:0] __delay_data_966_reinterpretcast_614;
  reg [1-1:0] __delay_data_967_pointer_630;
  reg signed [32-1:0] __delay_data_968_reinterpretcast_615;
  reg [1-1:0] __delay_data_969_pointer_632;
  reg signed [32-1:0] __delay_data_970_reinterpretcast_616;
  reg [1-1:0] __delay_data_971_pointer_634;
  reg signed [32-1:0] __delay_data_972_reinterpretcast_617;
  reg [1-1:0] __delay_data_973__variable_281;
  reg [10-1:0] __delay_data_998__variable_276;
  reg signed [32-1:0] __delay_data_1011_cond_297;
  reg signed [32-1:0] __delay_data_1030_cond_304;
  reg [1-1:0] __delay_data_1069_eq_873;
  wire signed [32-1:0] _cond_data_341;
  assign _cond_data_341 = (_eq_data_339)? __delay_data_946__variable_332 : 1'sd0;
  wire signed [32-1:0] _cond_data_345;
  assign _cond_data_345 = (_eq_data_343)? __delay_data_947__variable_331 : _cond_data_341;
  wire signed [32-1:0] _cond_data_348;
  assign _cond_data_348 = (_eq_data_346)? __delay_data_948__variable_330 : _cond_data_345;
  wire signed [32-1:0] _cond_data_351;
  assign _cond_data_351 = (_eq_data_349)? __delay_data_948__variable_330 : 1'sd0;
  wire signed [32-1:0] _cond_data_355;
  assign _cond_data_355 = (_eq_data_353)? __delay_data_946__variable_332 : _cond_data_351;
  wire signed [32-1:0] _cond_data_358;
  assign _cond_data_358 = (_eq_data_356)? __delay_data_947__variable_331 : _cond_data_355;
  wire signed [32-1:0] _cond_data_361;
  assign _cond_data_361 = (_eq_data_359)? __delay_data_947__variable_331 : 1'sd0;
  wire signed [32-1:0] _cond_data_365;
  assign _cond_data_365 = (_eq_data_363)? __delay_data_948__variable_330 : _cond_data_361;
  wire signed [32-1:0] _cond_data_368;
  assign _cond_data_368 = (_eq_data_366)? __delay_data_946__variable_332 : _cond_data_365;
  wire signed [32-1:0] _cond_data_371;
  assign _cond_data_371 = (_eq_data_369)? __delay_data_949__variable_335 : 1'sd0;
  wire signed [32-1:0] _cond_data_375;
  assign _cond_data_375 = (_eq_data_373)? __delay_data_950__variable_334 : _cond_data_371;
  wire signed [32-1:0] _cond_data_378;
  assign _cond_data_378 = (_eq_data_376)? __delay_data_951__variable_333 : _cond_data_375;
  wire signed [32-1:0] _cond_data_381;
  assign _cond_data_381 = (_eq_data_379)? __delay_data_951__variable_333 : 1'sd0;
  wire signed [32-1:0] _cond_data_385;
  assign _cond_data_385 = (_eq_data_383)? __delay_data_949__variable_335 : _cond_data_381;
  wire signed [32-1:0] _cond_data_388;
  assign _cond_data_388 = (_eq_data_386)? __delay_data_950__variable_334 : _cond_data_385;
  wire signed [32-1:0] _cond_data_391;
  assign _cond_data_391 = (_eq_data_389)? __delay_data_950__variable_334 : 1'sd0;
  wire signed [32-1:0] _cond_data_395;
  assign _cond_data_395 = (_eq_data_393)? __delay_data_951__variable_333 : _cond_data_391;
  wire signed [32-1:0] _cond_data_398;
  assign _cond_data_398 = (_eq_data_396)? __delay_data_949__variable_335 : _cond_data_395;
  wire signed [32-1:0] _cond_data_401;
  assign _cond_data_401 = (_eq_data_399)? __delay_data_952__variable_338 : 1'sd0;
  wire signed [32-1:0] _cond_data_405;
  assign _cond_data_405 = (_eq_data_403)? __delay_data_953__variable_337 : _cond_data_401;
  wire signed [32-1:0] _cond_data_408;
  assign _cond_data_408 = (_eq_data_406)? __delay_data_954__variable_336 : _cond_data_405;
  wire signed [32-1:0] _cond_data_411;
  assign _cond_data_411 = (_eq_data_409)? __delay_data_954__variable_336 : 1'sd0;
  wire signed [32-1:0] _cond_data_415;
  assign _cond_data_415 = (_eq_data_413)? __delay_data_952__variable_338 : _cond_data_411;
  wire signed [32-1:0] _cond_data_418;
  assign _cond_data_418 = (_eq_data_416)? __delay_data_953__variable_337 : _cond_data_415;
  wire signed [32-1:0] _cond_data_421;
  assign _cond_data_421 = (_eq_data_419)? __delay_data_953__variable_337 : 1'sd0;
  wire signed [32-1:0] _cond_data_425;
  assign _cond_data_425 = (_eq_data_423)? __delay_data_954__variable_336 : _cond_data_421;
  wire signed [32-1:0] _cond_data_428;
  assign _cond_data_428 = (_eq_data_426)? __delay_data_952__variable_338 : _cond_data_425;
  wire signed [32-1:0] _cond_data_431;
  assign _cond_data_431 = (_eq_data_429)? _cond_data_408 : 1'sd0;
  wire signed [32-1:0] _cond_data_435;
  assign _cond_data_435 = (_eq_data_433)? _cond_data_378 : _cond_data_431;
  wire signed [32-1:0] _cond_data_438;
  assign _cond_data_438 = (_eq_data_436)? _cond_data_348 : _cond_data_435;
  wire signed [32-1:0] _cond_data_441;
  assign _cond_data_441 = (_eq_data_439)? _cond_data_348 : 1'sd0;
  wire signed [32-1:0] _cond_data_445;
  assign _cond_data_445 = (_eq_data_443)? _cond_data_408 : _cond_data_441;
  wire signed [32-1:0] _cond_data_448;
  assign _cond_data_448 = (_eq_data_446)? _cond_data_378 : _cond_data_445;
  wire signed [32-1:0] _cond_data_451;
  assign _cond_data_451 = (_eq_data_449)? _cond_data_378 : 1'sd0;
  wire signed [32-1:0] _cond_data_455;
  assign _cond_data_455 = (_eq_data_453)? _cond_data_348 : _cond_data_451;
  wire signed [32-1:0] _cond_data_458;
  assign _cond_data_458 = (_eq_data_456)? _cond_data_408 : _cond_data_455;
  wire signed [32-1:0] _cond_data_461;
  assign _cond_data_461 = (_eq_data_459)? _cond_data_418 : 1'sd0;
  wire signed [32-1:0] _cond_data_465;
  assign _cond_data_465 = (_eq_data_463)? _cond_data_388 : _cond_data_461;
  wire signed [32-1:0] _cond_data_468;
  assign _cond_data_468 = (_eq_data_466)? _cond_data_358 : _cond_data_465;
  wire signed [32-1:0] _cond_data_471;
  assign _cond_data_471 = (_eq_data_469)? _cond_data_358 : 1'sd0;
  wire signed [32-1:0] _cond_data_475;
  assign _cond_data_475 = (_eq_data_473)? _cond_data_418 : _cond_data_471;
  wire signed [32-1:0] _cond_data_478;
  assign _cond_data_478 = (_eq_data_476)? _cond_data_388 : _cond_data_475;
  wire signed [32-1:0] _cond_data_481;
  assign _cond_data_481 = (_eq_data_479)? _cond_data_388 : 1'sd0;
  wire signed [32-1:0] _cond_data_485;
  assign _cond_data_485 = (_eq_data_483)? _cond_data_358 : _cond_data_481;
  wire signed [32-1:0] _cond_data_488;
  assign _cond_data_488 = (_eq_data_486)? _cond_data_418 : _cond_data_485;
  wire signed [32-1:0] _cond_data_491;
  assign _cond_data_491 = (_eq_data_489)? _cond_data_428 : 1'sd0;
  wire signed [32-1:0] _cond_data_495;
  assign _cond_data_495 = (_eq_data_493)? _cond_data_398 : _cond_data_491;
  wire signed [32-1:0] _cond_data_498;
  assign _cond_data_498 = (_eq_data_496)? _cond_data_368 : _cond_data_495;
  wire signed [32-1:0] _cond_data_501;
  assign _cond_data_501 = (_eq_data_499)? _cond_data_368 : 1'sd0;
  wire signed [32-1:0] _cond_data_505;
  assign _cond_data_505 = (_eq_data_503)? _cond_data_428 : _cond_data_501;
  wire signed [32-1:0] _cond_data_508;
  assign _cond_data_508 = (_eq_data_506)? _cond_data_398 : _cond_data_505;
  wire signed [32-1:0] _cond_data_511;
  assign _cond_data_511 = (_eq_data_509)? _cond_data_398 : 1'sd0;
  wire signed [32-1:0] _cond_data_515;
  assign _cond_data_515 = (_eq_data_513)? _cond_data_368 : _cond_data_511;
  wire signed [32-1:0] _cond_data_518;
  assign _cond_data_518 = (_eq_data_516)? _cond_data_428 : _cond_data_515;
  wire signed [32-1:0] _reinterpretcast_src_555;
  assign _reinterpretcast_src_555 = _cond_data_438;
  wire signed [32-1:0] _reinterpretcast_data_555;
  assign _reinterpretcast_data_555 = _reinterpretcast_src_555;
  wire signed [32-1:0] _reinterpretcast_src_556;
  assign _reinterpretcast_src_556 = _cond_data_468;
  wire signed [32-1:0] _reinterpretcast_data_556;
  assign _reinterpretcast_data_556 = _reinterpretcast_src_556;
  wire signed [32-1:0] _reinterpretcast_src_557;
  assign _reinterpretcast_src_557 = _cond_data_498;
  wire signed [32-1:0] _reinterpretcast_data_557;
  assign _reinterpretcast_data_557 = _reinterpretcast_src_557;
  wire signed [32-1:0] _reinterpretcast_src_558;
  assign _reinterpretcast_src_558 = _cond_data_448;
  wire signed [32-1:0] _reinterpretcast_data_558;
  assign _reinterpretcast_data_558 = _reinterpretcast_src_558;
  wire signed [32-1:0] _reinterpretcast_src_559;
  assign _reinterpretcast_src_559 = _cond_data_478;
  wire signed [32-1:0] _reinterpretcast_data_559;
  assign _reinterpretcast_data_559 = _reinterpretcast_src_559;
  wire signed [32-1:0] _reinterpretcast_src_560;
  assign _reinterpretcast_src_560 = _cond_data_508;
  wire signed [32-1:0] _reinterpretcast_data_560;
  assign _reinterpretcast_data_560 = _reinterpretcast_src_560;
  wire signed [32-1:0] _reinterpretcast_src_561;
  assign _reinterpretcast_src_561 = _cond_data_458;
  wire signed [32-1:0] _reinterpretcast_data_561;
  assign _reinterpretcast_data_561 = _reinterpretcast_src_561;
  wire signed [32-1:0] _reinterpretcast_src_562;
  assign _reinterpretcast_src_562 = _cond_data_488;
  wire signed [32-1:0] _reinterpretcast_data_562;
  assign _reinterpretcast_data_562 = _reinterpretcast_src_562;
  wire signed [32-1:0] _reinterpretcast_src_563;
  assign _reinterpretcast_src_563 = _cond_data_518;
  wire signed [32-1:0] _reinterpretcast_data_563;
  assign _reinterpretcast_data_563 = _reinterpretcast_src_563;
  wire signed [32-1:0] _cond_data_637;
  assign _cond_data_637 = (__delay_data_955_pointer_618)? 1'sd0 : _reinterpretcast_data_555;
  wire signed [32-1:0] _cond_data_639;
  assign _cond_data_639 = (__delay_data_957_pointer_620)? 1'sd0 : _reinterpretcast_data_556;
  wire signed [32-1:0] _cond_data_641;
  assign _cond_data_641 = (__delay_data_959_pointer_622)? 1'sd0 : _reinterpretcast_data_557;
  wire signed [32-1:0] _cond_data_643;
  assign _cond_data_643 = (__delay_data_961_pointer_624)? 1'sd0 : _reinterpretcast_data_558;
  wire signed [32-1:0] _cond_data_645;
  assign _cond_data_645 = (__delay_data_963_pointer_626)? 1'sd0 : _reinterpretcast_data_559;
  wire signed [32-1:0] _cond_data_647;
  assign _cond_data_647 = (__delay_data_965_pointer_628)? 1'sd0 : _reinterpretcast_data_560;
  wire signed [32-1:0] _cond_data_649;
  assign _cond_data_649 = (__delay_data_967_pointer_630)? 1'sd0 : _reinterpretcast_data_561;
  wire signed [32-1:0] _cond_data_651;
  assign _cond_data_651 = (__delay_data_969_pointer_632)? 1'sd0 : _reinterpretcast_data_562;
  wire signed [32-1:0] _cond_data_653;
  assign _cond_data_653 = (__delay_data_971_pointer_634)? 1'sd0 : _reinterpretcast_data_563;
  reg signed [32-1:0] __variable_wdata_80;
  assign mul_4_x_data = __variable_wdata_80;
  reg signed [32-1:0] __variable_wdata_81;
  assign mul_4_y_data = __variable_wdata_81;
  reg [6-1:0] __variable_wdata_82;
  assign mul_4_rshift_data = __variable_wdata_82;
  assign _mul_4_is_root = ((_stream_conv2d_25_busy)? 0 : 1) && 1;
  assign _mul_4_stream_oready = ((_stream_conv2d_25_busy)? _stream_conv2d_25_stream_oready : 1) && _mul_4_stream_internal_oready;
  reg signed [32-1:0] __variable_wdata_101;
  assign mul_5_x_data = __variable_wdata_101;
  reg signed [32-1:0] __variable_wdata_102;
  assign mul_5_y_data = __variable_wdata_102;
  reg [6-1:0] __variable_wdata_103;
  assign mul_5_rshift_data = __variable_wdata_103;
  assign _mul_5_is_root = ((_stream_conv2d_25_busy)? 0 : 1) && 1;
  assign _mul_5_stream_oready = ((_stream_conv2d_25_busy)? _stream_conv2d_25_stream_oready : 1) && _mul_5_stream_internal_oready;
  reg signed [32-1:0] __variable_wdata_122;
  assign mul_6_x_data = __variable_wdata_122;
  reg signed [32-1:0] __variable_wdata_123;
  assign mul_6_y_data = __variable_wdata_123;
  reg [6-1:0] __variable_wdata_124;
  assign mul_6_rshift_data = __variable_wdata_124;
  assign _mul_6_is_root = ((_stream_conv2d_25_busy)? 0 : 1) && 1;
  assign _mul_6_stream_oready = ((_stream_conv2d_25_busy)? _stream_conv2d_25_stream_oready : 1) && _mul_6_stream_internal_oready;
  reg signed [32-1:0] __variable_wdata_143;
  assign mul_7_x_data = __variable_wdata_143;
  reg signed [32-1:0] __variable_wdata_144;
  assign mul_7_y_data = __variable_wdata_144;
  reg [6-1:0] __variable_wdata_145;
  assign mul_7_rshift_data = __variable_wdata_145;
  assign _mul_7_is_root = ((_stream_conv2d_25_busy)? 0 : 1) && 1;
  assign _mul_7_stream_oready = ((_stream_conv2d_25_busy)? _stream_conv2d_25_stream_oready : 1) && _mul_7_stream_internal_oready;
  reg signed [32-1:0] __variable_wdata_164;
  assign mul_8_x_data = __variable_wdata_164;
  reg signed [32-1:0] __variable_wdata_165;
  assign mul_8_y_data = __variable_wdata_165;
  reg [6-1:0] __variable_wdata_166;
  assign mul_8_rshift_data = __variable_wdata_166;
  assign _mul_8_is_root = ((_stream_conv2d_25_busy)? 0 : 1) && 1;
  assign _mul_8_stream_oready = ((_stream_conv2d_25_busy)? _stream_conv2d_25_stream_oready : 1) && _mul_8_stream_internal_oready;
  reg signed [32-1:0] __variable_wdata_185;
  assign mul_9_x_data = __variable_wdata_185;
  reg signed [32-1:0] __variable_wdata_186;
  assign mul_9_y_data = __variable_wdata_186;
  reg [6-1:0] __variable_wdata_187;
  assign mul_9_rshift_data = __variable_wdata_187;
  assign _mul_9_is_root = ((_stream_conv2d_25_busy)? 0 : 1) && 1;
  assign _mul_9_stream_oready = ((_stream_conv2d_25_busy)? _stream_conv2d_25_stream_oready : 1) && _mul_9_stream_internal_oready;
  reg signed [32-1:0] __variable_wdata_206;
  assign mul_10_x_data = __variable_wdata_206;
  reg signed [32-1:0] __variable_wdata_207;
  assign mul_10_y_data = __variable_wdata_207;
  reg [6-1:0] __variable_wdata_208;
  assign mul_10_rshift_data = __variable_wdata_208;
  assign _mul_10_is_root = ((_stream_conv2d_25_busy)? 0 : 1) && 1;
  assign _mul_10_stream_oready = ((_stream_conv2d_25_busy)? _stream_conv2d_25_stream_oready : 1) && _mul_10_stream_internal_oready;
  reg signed [32-1:0] __variable_wdata_227;
  assign mul_11_x_data = __variable_wdata_227;
  reg signed [32-1:0] __variable_wdata_228;
  assign mul_11_y_data = __variable_wdata_228;
  reg [6-1:0] __variable_wdata_229;
  assign mul_11_rshift_data = __variable_wdata_229;
  assign _mul_11_is_root = ((_stream_conv2d_25_busy)? 0 : 1) && 1;
  assign _mul_11_stream_oready = ((_stream_conv2d_25_busy)? _stream_conv2d_25_stream_oready : 1) && _mul_11_stream_internal_oready;
  reg signed [32-1:0] __variable_wdata_248;
  assign mul_12_x_data = __variable_wdata_248;
  reg signed [32-1:0] __variable_wdata_249;
  assign mul_12_y_data = __variable_wdata_249;
  reg [6-1:0] __variable_wdata_250;
  assign mul_12_rshift_data = __variable_wdata_250;
  assign _mul_12_is_root = ((_stream_conv2d_25_busy)? 0 : 1) && 1;
  assign _mul_12_stream_oready = ((_stream_conv2d_25_busy)? _stream_conv2d_25_stream_oready : 1) && _mul_12_stream_internal_oready;
  reg [1-1:0] __delay_data_974__delay_973__variable_281;
  reg [32-1:0] __delay_data_986_plus_839;
  reg [10-1:0] __delay_data_999__delay_998__variable_276;
  reg signed [32-1:0] __delay_data_1012__delay_1011_cond_297;
  reg signed [32-1:0] __delay_data_1031__delay_1030_cond_304;
  reg [32-1:0] __delay_data_1050_plus_858;
  reg [1-1:0] __delay_data_1070__delay_1069_eq_873;
  reg [1-1:0] __delay_data_975__delay_974__delay_973__variable_281;
  reg [32-1:0] __delay_data_987__delay_986_plus_839;
  reg [10-1:0] __delay_data_1000__delay_999__delay_998__variable_276;
  reg signed [32-1:0] __delay_data_1013__delay_1012__delay_1011_cond_297;
  reg signed [32-1:0] __delay_data_1032__delay_1031__delay_1030_cond_304;
  reg [32-1:0] __delay_data_1051__delay_1050_plus_858;
  reg [1-1:0] __delay_data_1071__delay_1070__delay_1069_eq_873;
  reg [1-1:0] __delay_data_976__delay_975__delay_974____variable_281;
  reg [32-1:0] __delay_data_988__delay_987__delay_986_plus_839;
  reg [10-1:0] __delay_data_1001__delay_1000__delay_999____variable_276;
  reg signed [32-1:0] __delay_data_1014__delay_1013__delay_1012__delay_1011_cond_297;
  reg signed [32-1:0] __delay_data_1033__delay_1032__delay_1031__delay_1030_cond_304;
  reg [32-1:0] __delay_data_1052__delay_1051__delay_1050_plus_858;
  reg [1-1:0] __delay_data_1072__delay_1071__delay_1070__delay_1069_eq_873;
  reg [1-1:0] __delay_data_977__delay_976__delay_975____variable_281;
  reg [32-1:0] __delay_data_989__delay_988__delay_987__delay_986_plus_839;
  reg [10-1:0] __delay_data_1002__delay_1001__delay_1000____variable_276;
  reg signed [32-1:0] __delay_data_1015__delay_1014__delay_1013__delay_1012___cond_297;
  reg signed [32-1:0] __delay_data_1034__delay_1033__delay_1032__delay_1031___cond_304;
  reg [32-1:0] __delay_data_1053__delay_1052__delay_1051__delay_1050_plus_858;
  reg [1-1:0] __delay_data_1073__delay_1072__delay_1071__delay_1070___eq_873;
  reg [1-1:0] __delay_data_978__delay_977__delay_976____variable_281;
  reg [32-1:0] __delay_data_990__delay_989__delay_988__delay_987___plus_839;
  reg [10-1:0] __delay_data_1003__delay_1002__delay_1001____variable_276;
  reg signed [32-1:0] __delay_data_1016__delay_1015__delay_1014__delay_1013___cond_297;
  reg signed [32-1:0] __delay_data_1035__delay_1034__delay_1033__delay_1032___cond_304;
  reg [32-1:0] __delay_data_1054__delay_1053__delay_1052__delay_1051___plus_858;
  reg [1-1:0] __delay_data_1074__delay_1073__delay_1072__delay_1071___eq_873;
  reg [1-1:0] __delay_data_979__delay_978__delay_977____variable_281;
  reg [32-1:0] __delay_data_991__delay_990__delay_989__delay_988___plus_839;
  reg [10-1:0] __delay_data_1004__delay_1003__delay_1002____variable_276;
  reg signed [32-1:0] __delay_data_1017__delay_1016__delay_1015__delay_1014___cond_297;
  reg signed [32-1:0] __delay_data_1036__delay_1035__delay_1034__delay_1033___cond_304;
  reg [32-1:0] __delay_data_1055__delay_1054__delay_1053__delay_1052___plus_858;
  reg [1-1:0] __delay_data_1075__delay_1074__delay_1073__delay_1072___eq_873;
  reg [1-1:0] __delay_data_980__delay_979__delay_978____variable_281;
  reg [32-1:0] __delay_data_992__delay_991__delay_990__delay_989___plus_839;
  reg [10-1:0] __delay_data_1005__delay_1004__delay_1003____variable_276;
  reg signed [32-1:0] __delay_data_1018__delay_1017__delay_1016__delay_1015___cond_297;
  reg signed [32-1:0] __delay_data_1037__delay_1036__delay_1035__delay_1034___cond_304;
  reg [32-1:0] __delay_data_1056__delay_1055__delay_1054__delay_1053___plus_858;
  reg [1-1:0] __delay_data_1076__delay_1075__delay_1074__delay_1073___eq_873;
  reg [1-1:0] __delay_data_981__delay_980__delay_979____variable_281;
  reg [32-1:0] __delay_data_993__delay_992__delay_991__delay_990___plus_839;
  reg [10-1:0] __delay_data_1006__delay_1005__delay_1004____variable_276;
  reg signed [32-1:0] __delay_data_1019__delay_1018__delay_1017__delay_1016___cond_297;
  reg signed [32-1:0] __delay_data_1038__delay_1037__delay_1036__delay_1035___cond_304;
  reg [32-1:0] __delay_data_1057__delay_1056__delay_1055__delay_1054___plus_858;
  reg [1-1:0] __delay_data_1077__delay_1076__delay_1075__delay_1074___eq_873;
  reg [1-1:0] __delay_data_982__delay_981__delay_980____variable_281;
  reg [32-1:0] __delay_data_994__delay_993__delay_992__delay_991___plus_839;
  reg [10-1:0] __delay_data_1007__delay_1006__delay_1005____variable_276;
  reg signed [32-1:0] __delay_data_1020__delay_1019__delay_1018__delay_1017___cond_297;
  reg signed [32-1:0] __delay_data_1039__delay_1038__delay_1037__delay_1036___cond_304;
  reg [32-1:0] __delay_data_1058__delay_1057__delay_1056__delay_1055___plus_858;
  reg [1-1:0] __delay_data_1078__delay_1077__delay_1076__delay_1075___eq_873;
  wire signed [64-1:0] __substreamoutput_data_672;
  assign __substreamoutput_data_672 = mul_4_z_data;
  wire signed [64-1:0] __substreamoutput_data_691;
  assign __substreamoutput_data_691 = mul_5_z_data;
  wire signed [64-1:0] __substreamoutput_data_710;
  assign __substreamoutput_data_710 = mul_6_z_data;
  wire signed [64-1:0] __substreamoutput_data_729;
  assign __substreamoutput_data_729 = mul_7_z_data;
  wire signed [64-1:0] __substreamoutput_data_748;
  assign __substreamoutput_data_748 = mul_8_z_data;
  wire signed [64-1:0] __substreamoutput_data_767;
  assign __substreamoutput_data_767 = mul_9_z_data;
  wire signed [64-1:0] __substreamoutput_data_786;
  assign __substreamoutput_data_786 = mul_10_z_data;
  wire signed [64-1:0] __substreamoutput_data_805;
  assign __substreamoutput_data_805 = mul_11_z_data;
  wire signed [64-1:0] __substreamoutput_data_824;
  assign __substreamoutput_data_824 = mul_12_z_data;
  reg signed [128-1:0] __variable_wdata_32;
  assign add_tree_2_var0_data = __variable_wdata_32;
  reg signed [128-1:0] __variable_wdata_33;
  assign add_tree_2_var1_data = __variable_wdata_33;
  reg signed [128-1:0] __variable_wdata_34;
  assign add_tree_2_var2_data = __variable_wdata_34;
  reg signed [128-1:0] __variable_wdata_35;
  assign add_tree_2_var3_data = __variable_wdata_35;
  reg signed [128-1:0] __variable_wdata_36;
  assign add_tree_2_var4_data = __variable_wdata_36;
  reg signed [128-1:0] __variable_wdata_37;
  assign add_tree_2_var5_data = __variable_wdata_37;
  reg signed [128-1:0] __variable_wdata_38;
  assign add_tree_2_var6_data = __variable_wdata_38;
  reg signed [128-1:0] __variable_wdata_39;
  assign add_tree_2_var7_data = __variable_wdata_39;
  reg signed [128-1:0] __variable_wdata_40;
  assign add_tree_2_var8_data = __variable_wdata_40;
  assign _add_tree_2_is_root = ((_stream_conv2d_25_busy)? 0 : 1) && 1;
  assign _add_tree_2_stream_oready = ((_stream_conv2d_25_busy)? _stream_conv2d_25_stream_oready : 1) && _add_tree_2_stream_internal_oready;
  reg [1-1:0] __delay_data_983__delay_982__delay_981____variable_281;
  reg [32-1:0] __delay_data_995__delay_994__delay_993__delay_992___plus_839;
  reg [10-1:0] __delay_data_1008__delay_1007__delay_1006____variable_276;
  reg signed [32-1:0] __delay_data_1021__delay_1020__delay_1019__delay_1018___cond_297;
  reg signed [32-1:0] __delay_data_1040__delay_1039__delay_1038__delay_1037___cond_304;
  reg [32-1:0] __delay_data_1059__delay_1058__delay_1057__delay_1056___plus_858;
  reg [1-1:0] __delay_data_1079__delay_1078__delay_1077__delay_1076___eq_873;
  reg [1-1:0] __delay_data_984__delay_983__delay_982____variable_281;
  reg [32-1:0] __delay_data_996__delay_995__delay_994__delay_993___plus_839;
  reg [10-1:0] __delay_data_1009__delay_1008__delay_1007____variable_276;
  reg signed [32-1:0] __delay_data_1022__delay_1021__delay_1020__delay_1019___cond_297;
  reg signed [32-1:0] __delay_data_1041__delay_1040__delay_1039__delay_1038___cond_304;
  reg [32-1:0] __delay_data_1060__delay_1059__delay_1058__delay_1057___plus_858;
  reg [1-1:0] __delay_data_1080__delay_1079__delay_1078__delay_1077___eq_873;
  reg [1-1:0] __delay_data_985__delay_984__delay_983____variable_281;
  reg [32-1:0] __delay_data_997__delay_996__delay_995__delay_994___plus_839;
  reg [10-1:0] __delay_data_1010__delay_1009__delay_1008____variable_276;
  reg signed [32-1:0] __delay_data_1023__delay_1022__delay_1021__delay_1020___cond_297;
  reg signed [32-1:0] __delay_data_1042__delay_1041__delay_1040__delay_1039___cond_304;
  reg [32-1:0] __delay_data_1061__delay_1060__delay_1059__delay_1058___plus_858;
  reg [1-1:0] __delay_data_1081__delay_1080__delay_1079__delay_1078___eq_873;
  wire signed [128-1:0] __substreamoutput_data_826;
  assign __substreamoutput_data_826 = add_tree_2_sum_data;
  reg [1-1:0] __variable_wdata_25;
  assign acc_1__reduce_reset_data = __variable_wdata_25;
  reg signed [128-1:0] __variable_wdata_10;
  assign acc_1_x_data = __variable_wdata_10;
  reg [8-1:0] __variable_wdata_11;
  assign acc_1_rshift_data = __variable_wdata_11;
  reg [32-1:0] __variable_wdata_12;
  assign acc_1_size_data = __variable_wdata_12;
  assign _acc_1_is_root = ((_stream_conv2d_25_busy)? 0 : 1) && 1;
  assign _acc_1_stream_oready = ((_stream_conv2d_25_busy)? _stream_conv2d_25_stream_oready : 1) && _acc_1_stream_internal_oready;
  reg signed [32-1:0] __delay_data_1024__delay_1023__delay_1022__delay_1021___cond_297;
  reg signed [32-1:0] __delay_data_1043__delay_1042__delay_1041__delay_1040___cond_304;
  reg [32-1:0] __delay_data_1062__delay_1061__delay_1060__delay_1059___plus_858;
  reg [1-1:0] __delay_data_1082__delay_1081__delay_1080__delay_1079___eq_873;
  reg signed [32-1:0] __delay_data_1025__delay_1024__delay_1023__delay_1022___cond_297;
  reg signed [32-1:0] __delay_data_1044__delay_1043__delay_1042__delay_1041___cond_304;
  reg [32-1:0] __delay_data_1063__delay_1062__delay_1061__delay_1060___plus_858;
  reg [1-1:0] __delay_data_1083__delay_1082__delay_1081__delay_1080___eq_873;
  reg signed [32-1:0] __delay_data_1026__delay_1025__delay_1024__delay_1023___cond_297;
  reg signed [32-1:0] __delay_data_1045__delay_1044__delay_1043__delay_1042___cond_304;
  reg [32-1:0] __delay_data_1064__delay_1063__delay_1062__delay_1061___plus_858;
  reg [1-1:0] __delay_data_1084__delay_1083__delay_1082__delay_1081___eq_873;
  reg signed [32-1:0] __delay_data_1027__delay_1026__delay_1025__delay_1024___cond_297;
  reg signed [32-1:0] __delay_data_1046__delay_1045__delay_1044__delay_1043___cond_304;
  reg [32-1:0] __delay_data_1065__delay_1064__delay_1063__delay_1062___plus_858;
  reg [1-1:0] __delay_data_1085__delay_1084__delay_1083__delay_1082___eq_873;
  reg signed [32-1:0] __delay_data_1028__delay_1027__delay_1026__delay_1025___cond_297;
  reg signed [32-1:0] __delay_data_1047__delay_1046__delay_1045__delay_1044___cond_304;
  reg [32-1:0] __delay_data_1066__delay_1065__delay_1064__delay_1063___plus_858;
  reg [1-1:0] __delay_data_1086__delay_1085__delay_1084__delay_1083___eq_873;
  reg signed [32-1:0] __delay_data_1029__delay_1028__delay_1027__delay_1026___cond_297;
  reg signed [32-1:0] __delay_data_1048__delay_1047__delay_1046__delay_1045___cond_304;
  reg [32-1:0] __delay_data_1067__delay_1066__delay_1065__delay_1064___plus_858;
  reg [1-1:0] __delay_data_1087__delay_1086__delay_1085__delay_1084___eq_873;
  wire signed [128-1:0] __substreamoutput_data_840;
  assign __substreamoutput_data_840 = acc_1_sum_data;
  wire [1-1:0] __substreamoutput_data_841;
  assign __substreamoutput_data_841 = acc_1_valid_data;
  reg signed [128-1:0] _plus_data_842;
  reg signed [32-1:0] __delay_data_1049__delay_1048__delay_1047__delay_1046___cond_304;
  reg [32-1:0] __delay_data_1068__delay_1067__delay_1066__delay_1065___plus_858;
  reg [1-1:0] __delay_data_1088__delay_1087__delay_1086__delay_1085___eq_873;
  reg [1-1:0] __delay_data_1108__substreamoutput_841;
  reg signed [128-1:0] __variable_wdata_46;
  assign mul_rshift_round_clip_3_x_data = __variable_wdata_46;
  reg signed [32-1:0] __variable_wdata_47;
  assign mul_rshift_round_clip_3_y_data = __variable_wdata_47;
  reg [8-1:0] __variable_wdata_48;
  assign mul_rshift_round_clip_3_rshift_data = __variable_wdata_48;
  assign _mul_rshift_round_clip_3_is_root = ((_stream_conv2d_25_busy)? 0 : 1) && 1;
  assign _mul_rshift_round_clip_3_stream_oready = ((_stream_conv2d_25_busy)? _stream_conv2d_25_stream_oready : 1) && _mul_rshift_round_clip_3_stream_internal_oready;
  assign _stream_conv2d_25_stream_internal_oready = ((_stream_conv2d_25_busy)? _mul_rshift_round_clip_3_stream_internal_oready : 1) && (((_stream_conv2d_25_busy)? _acc_1_stream_internal_oready : 1) && (((_stream_conv2d_25_busy)? _add_tree_2_stream_internal_oready : 1) && (((_stream_conv2d_25_busy)? _mul_12_stream_internal_oready : 1) && (((_stream_conv2d_25_busy)? _mul_11_stream_internal_oready : 1) && (((_stream_conv2d_25_busy)? _mul_10_stream_internal_oready : 1) && (((_stream_conv2d_25_busy)? _mul_9_stream_internal_oready : 1) && (((_stream_conv2d_25_busy)? _mul_8_stream_internal_oready : 1) && (((_stream_conv2d_25_busy)? _mul_7_stream_internal_oready : 1) && (((_stream_conv2d_25_busy)? _mul_6_stream_internal_oready : 1) && (((_stream_conv2d_25_busy)? _mul_5_stream_internal_oready : 1) && (((_stream_conv2d_25_busy)? _mul_4_stream_internal_oready : 1) && 1)))))))))));
  reg [1-1:0] __delay_data_1089__delay_1088__delay_1087__delay_1086___eq_873;
  reg [1-1:0] __delay_data_1109__delay_1108__substreamoutput_841;
  reg [1-1:0] __delay_data_1090__delay_1089__delay_1088__delay_1087___eq_873;
  reg [1-1:0] __delay_data_1110__delay_1109__delay_1108__substreamoutput_841;
  reg [1-1:0] __delay_data_1091__delay_1090__delay_1089__delay_1088___eq_873;
  reg [1-1:0] __delay_data_1111__delay_1110__delay_1109____substreamoutput_841;
  reg [1-1:0] __delay_data_1092__delay_1091__delay_1090__delay_1089___eq_873;
  reg [1-1:0] __delay_data_1112__delay_1111__delay_1110____substreamoutput_841;
  reg [1-1:0] __delay_data_1093__delay_1092__delay_1091__delay_1090___eq_873;
  reg [1-1:0] __delay_data_1113__delay_1112__delay_1111____substreamoutput_841;
  reg [1-1:0] __delay_data_1094__delay_1093__delay_1092__delay_1091___eq_873;
  reg [1-1:0] __delay_data_1114__delay_1113__delay_1112____substreamoutput_841;
  reg [1-1:0] __delay_data_1095__delay_1094__delay_1093__delay_1092___eq_873;
  reg [1-1:0] __delay_data_1115__delay_1114__delay_1113____substreamoutput_841;
  reg [1-1:0] __delay_data_1096__delay_1095__delay_1094__delay_1093___eq_873;
  reg [1-1:0] __delay_data_1116__delay_1115__delay_1114____substreamoutput_841;
  reg [1-1:0] __delay_data_1097__delay_1096__delay_1095__delay_1094___eq_873;
  reg [1-1:0] __delay_data_1117__delay_1116__delay_1115____substreamoutput_841;
  wire signed [32-1:0] __substreamoutput_data_859;
  assign __substreamoutput_data_859 = mul_rshift_round_clip_3_z_data;
  wire signed [61-1:0] _times_mul_odata_860;
  reg signed [61-1:0] _times_mul_odata_reg_860;
  wire signed [62-1:0] _times_data_860;
  assign _times_data_860 = _times_mul_odata_reg_860;
  wire _times_mul_update_860;
  assign _times_mul_update_860 = _stream_conv2d_25_stream_oready;

  multiplier_1
  _times_mul_860
  (
    .CLK(CLK),
    .update(_times_mul_update_860),
    .a(__substreamoutput_data_859),
    .b(29'sd214748368),
    .c(_times_mul_odata_860)
  );

  reg [1-1:0] _greaterthan_data_877;
  reg [1-1:0] __delay_data_1098__delay_1097__delay_1096__delay_1095___eq_873;
  reg signed [32-1:0] __delay_data_1104__substreamoutput_859;
  reg [1-1:0] __delay_data_1118__delay_1117__delay_1116____substreamoutput_841;
  reg [1-1:0] __delay_data_1099__delay_1098__delay_1097__delay_1096___eq_873;
  reg [1-1:0] __delay_data_1101_greaterthan_877;
  reg signed [32-1:0] __delay_data_1105__delay_1104__substreamoutput_859;
  reg [1-1:0] __delay_data_1119__delay_1118__delay_1117____substreamoutput_841;
  reg [1-1:0] __delay_data_1100__delay_1099__delay_1098__delay_1097___eq_873;
  reg [1-1:0] __delay_data_1102__delay_1101_greaterthan_877;
  reg signed [32-1:0] __delay_data_1106__delay_1105__delay_1104__substreamoutput_859;
  reg [1-1:0] __delay_data_1120__delay_1119__delay_1118____substreamoutput_841;
  wire [1-1:0] _pointer_data_862;
  assign _pointer_data_862 = _times_data_860[7'sd61];
  wire signed [2-1:0] _cond_data_866;
  assign _cond_data_866 = (_pointer_data_862)? -2'sd1 : 1'sd0;
  wire signed [63-1:0] _plus_data_867;
  assign _plus_data_867 = _times_data_860 + 32'sd1073741824;
  wire signed [63-1:0] _plus_data_869;
  assign _plus_data_869 = _plus_data_867 + _cond_data_866;
  wire signed [62-1:0] _sra_data_870;
  assign _sra_data_870 = _plus_data_869 >>> 6'sd31;
  reg signed [32-1:0] _cond_data_875;
  reg [1-1:0] __delay_data_1103__delay_1102__delay_1101_greaterthan_877;
  reg signed [32-1:0] __delay_data_1107__delay_1106__delay_1105____substreamoutput_859;
  reg [1-1:0] __delay_data_1121__delay_1120__delay_1119____substreamoutput_841;
  reg signed [32-1:0] _cond_data_878;
  reg [1-1:0] __delay_data_1122__delay_1121__delay_1120____substreamoutput_841;
  wire signed [32-1:0] _reinterpretcast_src_879;
  assign _reinterpretcast_src_879 = _cond_data_878;
  wire signed [32-1:0] _reinterpretcast_data_879;
  assign _reinterpretcast_data_879 = _reinterpretcast_src_879;
  wire signed [32-1:0] stream_conv2d_25_sink_50_data;
  assign stream_conv2d_25_sink_50_data = _reinterpretcast_data_879;
  wire [1-1:0] stream_conv2d_25_sink_51_data;
  assign stream_conv2d_25_sink_51_data = __delay_data_1122__delay_1121__delay_1120____substreamoutput_841;
  wire _set_flag_218;
  assign _set_flag_218 = conv2d_25_comp_fsm == 3;
  reg [10-1:0] __variable_wdata_276;
  assign stream_conv2d_25_parameter_0_data = __variable_wdata_276;
  wire _set_flag_219;
  assign _set_flag_219 = conv2d_25_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_277;
  assign stream_conv2d_25_parameter_1_data = __variable_wdata_277;
  wire _set_flag_220;
  assign _set_flag_220 = conv2d_25_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_278;
  assign stream_conv2d_25_parameter_2_data = __variable_wdata_278;
  wire _set_flag_221;
  assign _set_flag_221 = conv2d_25_comp_fsm == 3;
  reg [9-1:0] __variable_wdata_279;
  assign stream_conv2d_25_parameter_3_data = __variable_wdata_279;
  wire _set_flag_222;
  assign _set_flag_222 = conv2d_25_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_280;
  assign stream_conv2d_25_parameter_4_data = __variable_wdata_280;
  wire _set_flag_223;
  assign _set_flag_223 = conv2d_25_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_291;
  assign stream_conv2d_25_parameter_6_data = __variable_wdata_291;
  reg [32-1:0] _source_stream_conv2d_25_source_7_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_7_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_7_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_7_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_7_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_7_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_7_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_7_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_7_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_7_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_7_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_7_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_7_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_7_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_7_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_7_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_7_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_7_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_7_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_7_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_7_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_7_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_7_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_7_pat_stride_buf_3;
  wire _set_flag_224;
  assign _set_flag_224 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l4096_id0_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_7_source_ram_renable && (_stream_conv2d_25_source_7_source_sel == 1))? _stream_conv2d_25_source_7_source_ram_raddr : 'hx;
  assign ram_w32_l4096_id0_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_7_source_ram_renable && (_stream_conv2d_25_source_7_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_225 = 1;
  wire [_tmp_225-1:0] _tmp_226;
  assign _tmp_226 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_7_source_ram_renable && (_stream_conv2d_25_source_7_source_sel == 1);
  reg [_tmp_225-1:0] __tmp_226_1;
  assign _stream_conv2d_25_source_7_source_ram_rdata = (_stream_conv2d_25_source_7_source_sel == 1)? ram_w32_l4096_id0_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_292;
  assign stream_conv2d_25_source_7_data = __variable_wdata_292;
  reg [32-1:0] _stream_conv2d_25_source_7_source_pat_fsm_0;
  localparam _stream_conv2d_25_source_7_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_7_source_pat_all_offset;
  assign _stream_conv2d_25_source_7_source_pat_all_offset = _stream_conv2d_25_source_7_source_offset_buf + _source_stream_conv2d_25_source_7_pat_cur_offset_0 + _source_stream_conv2d_25_source_7_pat_cur_offset_1 + _source_stream_conv2d_25_source_7_pat_cur_offset_2 + _source_stream_conv2d_25_source_7_pat_cur_offset_3;
  wire _set_flag_227;
  assign _set_flag_227 = conv2d_25_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_298;
  assign stream_conv2d_25_parameter_8_data = __variable_wdata_298;
  reg [32-1:0] _source_stream_conv2d_25_source_9_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_9_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_9_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_9_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_9_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_9_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_9_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_9_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_9_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_9_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_9_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_9_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_9_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_9_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_9_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_9_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_9_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_9_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_9_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_9_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_9_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_9_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_9_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_9_pat_stride_buf_3;
  wire _set_flag_228;
  assign _set_flag_228 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l1024_id0_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_9_source_ram_renable && (_stream_conv2d_25_source_9_source_sel == 2))? _stream_conv2d_25_source_9_source_ram_raddr : 'hx;
  assign ram_w32_l1024_id0_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_9_source_ram_renable && (_stream_conv2d_25_source_9_source_sel == 2))? 1'd1 : 0;
  localparam _tmp_229 = 1;
  wire [_tmp_229-1:0] _tmp_230;
  assign _tmp_230 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_9_source_ram_renable && (_stream_conv2d_25_source_9_source_sel == 2);
  reg [_tmp_229-1:0] __tmp_230_1;
  assign _stream_conv2d_25_source_9_source_ram_rdata = (_stream_conv2d_25_source_9_source_sel == 2)? ram_w32_l1024_id0_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_299;
  assign stream_conv2d_25_source_9_data = __variable_wdata_299;
  reg [32-1:0] _stream_conv2d_25_source_9_source_pat_fsm_1;
  localparam _stream_conv2d_25_source_9_source_pat_fsm_1_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_9_source_pat_all_offset;
  assign _stream_conv2d_25_source_9_source_pat_all_offset = _stream_conv2d_25_source_9_source_offset_buf + _source_stream_conv2d_25_source_9_pat_cur_offset_0 + _source_stream_conv2d_25_source_9_pat_cur_offset_1 + _source_stream_conv2d_25_source_9_pat_cur_offset_2 + _source_stream_conv2d_25_source_9_pat_cur_offset_3;
  wire _set_flag_231;
  assign _set_flag_231 = conv2d_25_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_305;
  assign stream_conv2d_25_parameter_10_data = __variable_wdata_305;
  wire _set_flag_232;
  assign _set_flag_232 = conv2d_25_comp_fsm == 3;
  reg [32-1:0] __variable_wdata_306;
  assign stream_conv2d_25_source_11_data = __variable_wdata_306;
  wire _set_flag_233;
  assign _set_flag_233 = conv2d_25_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_312;
  assign stream_conv2d_25_parameter_12_data = __variable_wdata_312;
  wire _set_flag_234;
  assign _set_flag_234 = conv2d_25_comp_fsm == 3;
  reg [32-1:0] __variable_wdata_313;
  assign stream_conv2d_25_source_13_data = __variable_wdata_313;
  wire _set_flag_235;
  assign _set_flag_235 = conv2d_25_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_319;
  assign stream_conv2d_25_parameter_14_data = __variable_wdata_319;
  wire _set_flag_236;
  assign _set_flag_236 = conv2d_25_comp_fsm == 3;
  reg [32-1:0] __variable_wdata_320;
  assign stream_conv2d_25_source_15_data = __variable_wdata_320;
  wire _set_flag_237;
  assign _set_flag_237 = conv2d_25_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_326;
  assign stream_conv2d_25_parameter_16_data = __variable_wdata_326;
  wire _set_flag_238;
  assign _set_flag_238 = conv2d_25_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_327;
  assign stream_conv2d_25_parameter_17_data = __variable_wdata_327;
  wire _set_flag_239;
  assign _set_flag_239 = conv2d_25_comp_fsm == 3;
  reg [5-1:0] __variable_wdata_328;
  assign stream_conv2d_25_parameter_18_data = __variable_wdata_328;
  wire _set_flag_240;
  assign _set_flag_240 = conv2d_25_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_329;
  assign stream_conv2d_25_parameter_19_data = __variable_wdata_329;
  reg [32-1:0] _source_stream_conv2d_25_source_20_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_20_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_20_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_20_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_20_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_20_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_20_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_20_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_20_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_20_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_20_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_20_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_20_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_20_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_20_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_20_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_20_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_20_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_20_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_20_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_20_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_20_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_20_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_20_pat_stride_buf_3;
  wire _set_flag_241;
  assign _set_flag_241 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l4096_id1_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_20_source_ram_renable && (_stream_conv2d_25_source_20_source_sel == 3))? _stream_conv2d_25_source_20_source_ram_raddr : 'hx;
  assign ram_w32_l4096_id1_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_20_source_ram_renable && (_stream_conv2d_25_source_20_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_242 = 1;
  wire [_tmp_242-1:0] _tmp_243;
  assign _tmp_243 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_20_source_ram_renable && (_stream_conv2d_25_source_20_source_sel == 3);
  reg [_tmp_242-1:0] __tmp_243_1;
  assign _stream_conv2d_25_source_20_source_ram_rdata = (_stream_conv2d_25_source_20_source_sel == 3)? ram_w32_l4096_id1_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_330;
  assign stream_conv2d_25_source_20_data = __variable_wdata_330;
  reg [32-1:0] _stream_conv2d_25_source_20_source_pat_fsm_2;
  localparam _stream_conv2d_25_source_20_source_pat_fsm_2_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_20_source_pat_all_offset;
  assign _stream_conv2d_25_source_20_source_pat_all_offset = _stream_conv2d_25_source_20_source_offset_buf + _source_stream_conv2d_25_source_20_pat_cur_offset_0 + _source_stream_conv2d_25_source_20_pat_cur_offset_1 + _source_stream_conv2d_25_source_20_pat_cur_offset_2 + _source_stream_conv2d_25_source_20_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_25_source_21_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_21_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_21_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_21_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_21_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_21_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_21_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_21_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_21_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_21_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_21_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_21_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_21_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_21_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_21_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_21_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_21_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_21_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_21_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_21_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_21_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_21_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_21_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_21_pat_stride_buf_3;
  wire _set_flag_244;
  assign _set_flag_244 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l4096_id2_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_21_source_ram_renable && (_stream_conv2d_25_source_21_source_sel == 4))? _stream_conv2d_25_source_21_source_ram_raddr : 'hx;
  assign ram_w32_l4096_id2_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_21_source_ram_renable && (_stream_conv2d_25_source_21_source_sel == 4))? 1'd1 : 0;
  localparam _tmp_245 = 1;
  wire [_tmp_245-1:0] _tmp_246;
  assign _tmp_246 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_21_source_ram_renable && (_stream_conv2d_25_source_21_source_sel == 4);
  reg [_tmp_245-1:0] __tmp_246_1;
  assign _stream_conv2d_25_source_21_source_ram_rdata = (_stream_conv2d_25_source_21_source_sel == 4)? ram_w32_l4096_id2_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_331;
  assign stream_conv2d_25_source_21_data = __variable_wdata_331;
  reg [32-1:0] _stream_conv2d_25_source_21_source_pat_fsm_3;
  localparam _stream_conv2d_25_source_21_source_pat_fsm_3_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_21_source_pat_all_offset;
  assign _stream_conv2d_25_source_21_source_pat_all_offset = _stream_conv2d_25_source_21_source_offset_buf + _source_stream_conv2d_25_source_21_pat_cur_offset_0 + _source_stream_conv2d_25_source_21_pat_cur_offset_1 + _source_stream_conv2d_25_source_21_pat_cur_offset_2 + _source_stream_conv2d_25_source_21_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_25_source_22_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_22_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_22_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_22_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_22_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_22_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_22_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_22_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_22_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_22_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_22_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_22_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_22_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_22_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_22_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_22_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_22_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_22_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_22_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_22_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_22_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_22_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_22_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_22_pat_stride_buf_3;
  wire _set_flag_247;
  assign _set_flag_247 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l4096_id3_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_22_source_ram_renable && (_stream_conv2d_25_source_22_source_sel == 5))? _stream_conv2d_25_source_22_source_ram_raddr : 'hx;
  assign ram_w32_l4096_id3_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_22_source_ram_renable && (_stream_conv2d_25_source_22_source_sel == 5))? 1'd1 : 0;
  localparam _tmp_248 = 1;
  wire [_tmp_248-1:0] _tmp_249;
  assign _tmp_249 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_22_source_ram_renable && (_stream_conv2d_25_source_22_source_sel == 5);
  reg [_tmp_248-1:0] __tmp_249_1;
  assign _stream_conv2d_25_source_22_source_ram_rdata = (_stream_conv2d_25_source_22_source_sel == 5)? ram_w32_l4096_id3_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_332;
  assign stream_conv2d_25_source_22_data = __variable_wdata_332;
  reg [32-1:0] _stream_conv2d_25_source_22_source_pat_fsm_4;
  localparam _stream_conv2d_25_source_22_source_pat_fsm_4_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_22_source_pat_all_offset;
  assign _stream_conv2d_25_source_22_source_pat_all_offset = _stream_conv2d_25_source_22_source_offset_buf + _source_stream_conv2d_25_source_22_pat_cur_offset_0 + _source_stream_conv2d_25_source_22_pat_cur_offset_1 + _source_stream_conv2d_25_source_22_pat_cur_offset_2 + _source_stream_conv2d_25_source_22_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_25_source_23_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_23_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_23_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_23_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_23_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_23_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_23_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_23_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_23_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_23_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_23_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_23_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_23_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_23_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_23_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_23_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_23_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_23_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_23_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_23_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_23_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_23_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_23_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_23_pat_stride_buf_3;
  wire _set_flag_250;
  assign _set_flag_250 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l4096_id4_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_23_source_ram_renable && (_stream_conv2d_25_source_23_source_sel == 6))? _stream_conv2d_25_source_23_source_ram_raddr : 'hx;
  assign ram_w32_l4096_id4_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_23_source_ram_renable && (_stream_conv2d_25_source_23_source_sel == 6))? 1'd1 : 0;
  localparam _tmp_251 = 1;
  wire [_tmp_251-1:0] _tmp_252;
  assign _tmp_252 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_23_source_ram_renable && (_stream_conv2d_25_source_23_source_sel == 6);
  reg [_tmp_251-1:0] __tmp_252_1;
  assign _stream_conv2d_25_source_23_source_ram_rdata = (_stream_conv2d_25_source_23_source_sel == 6)? ram_w32_l4096_id4_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_333;
  assign stream_conv2d_25_source_23_data = __variable_wdata_333;
  reg [32-1:0] _stream_conv2d_25_source_23_source_pat_fsm_5;
  localparam _stream_conv2d_25_source_23_source_pat_fsm_5_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_23_source_pat_all_offset;
  assign _stream_conv2d_25_source_23_source_pat_all_offset = _stream_conv2d_25_source_23_source_offset_buf + _source_stream_conv2d_25_source_23_pat_cur_offset_0 + _source_stream_conv2d_25_source_23_pat_cur_offset_1 + _source_stream_conv2d_25_source_23_pat_cur_offset_2 + _source_stream_conv2d_25_source_23_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_25_source_24_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_24_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_24_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_24_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_24_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_24_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_24_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_24_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_24_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_24_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_24_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_24_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_24_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_24_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_24_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_24_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_24_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_24_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_24_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_24_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_24_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_24_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_24_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_24_pat_stride_buf_3;
  wire _set_flag_253;
  assign _set_flag_253 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l4096_id5_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_24_source_ram_renable && (_stream_conv2d_25_source_24_source_sel == 7))? _stream_conv2d_25_source_24_source_ram_raddr : 'hx;
  assign ram_w32_l4096_id5_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_24_source_ram_renable && (_stream_conv2d_25_source_24_source_sel == 7))? 1'd1 : 0;
  localparam _tmp_254 = 1;
  wire [_tmp_254-1:0] _tmp_255;
  assign _tmp_255 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_24_source_ram_renable && (_stream_conv2d_25_source_24_source_sel == 7);
  reg [_tmp_254-1:0] __tmp_255_1;
  assign _stream_conv2d_25_source_24_source_ram_rdata = (_stream_conv2d_25_source_24_source_sel == 7)? ram_w32_l4096_id5_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_334;
  assign stream_conv2d_25_source_24_data = __variable_wdata_334;
  reg [32-1:0] _stream_conv2d_25_source_24_source_pat_fsm_6;
  localparam _stream_conv2d_25_source_24_source_pat_fsm_6_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_24_source_pat_all_offset;
  assign _stream_conv2d_25_source_24_source_pat_all_offset = _stream_conv2d_25_source_24_source_offset_buf + _source_stream_conv2d_25_source_24_pat_cur_offset_0 + _source_stream_conv2d_25_source_24_pat_cur_offset_1 + _source_stream_conv2d_25_source_24_pat_cur_offset_2 + _source_stream_conv2d_25_source_24_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_25_source_25_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_25_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_25_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_25_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_25_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_25_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_25_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_25_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_25_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_25_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_25_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_25_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_25_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_25_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_25_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_25_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_25_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_25_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_25_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_25_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_25_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_25_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_25_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_25_pat_stride_buf_3;
  wire _set_flag_256;
  assign _set_flag_256 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l4096_id6_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_25_source_ram_renable && (_stream_conv2d_25_source_25_source_sel == 8))? _stream_conv2d_25_source_25_source_ram_raddr : 'hx;
  assign ram_w32_l4096_id6_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_25_source_ram_renable && (_stream_conv2d_25_source_25_source_sel == 8))? 1'd1 : 0;
  localparam _tmp_257 = 1;
  wire [_tmp_257-1:0] _tmp_258;
  assign _tmp_258 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_25_source_ram_renable && (_stream_conv2d_25_source_25_source_sel == 8);
  reg [_tmp_257-1:0] __tmp_258_1;
  assign _stream_conv2d_25_source_25_source_ram_rdata = (_stream_conv2d_25_source_25_source_sel == 8)? ram_w32_l4096_id6_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_335;
  assign stream_conv2d_25_source_25_data = __variable_wdata_335;
  reg [32-1:0] _stream_conv2d_25_source_25_source_pat_fsm_7;
  localparam _stream_conv2d_25_source_25_source_pat_fsm_7_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_25_source_pat_all_offset;
  assign _stream_conv2d_25_source_25_source_pat_all_offset = _stream_conv2d_25_source_25_source_offset_buf + _source_stream_conv2d_25_source_25_pat_cur_offset_0 + _source_stream_conv2d_25_source_25_pat_cur_offset_1 + _source_stream_conv2d_25_source_25_pat_cur_offset_2 + _source_stream_conv2d_25_source_25_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_25_source_26_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_26_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_26_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_26_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_26_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_26_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_26_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_26_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_26_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_26_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_26_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_26_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_26_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_26_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_26_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_26_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_26_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_26_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_26_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_26_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_26_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_26_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_26_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_26_pat_stride_buf_3;
  wire _set_flag_259;
  assign _set_flag_259 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l4096_id7_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_26_source_ram_renable && (_stream_conv2d_25_source_26_source_sel == 9))? _stream_conv2d_25_source_26_source_ram_raddr : 'hx;
  assign ram_w32_l4096_id7_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_26_source_ram_renable && (_stream_conv2d_25_source_26_source_sel == 9))? 1'd1 : 0;
  localparam _tmp_260 = 1;
  wire [_tmp_260-1:0] _tmp_261;
  assign _tmp_261 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_26_source_ram_renable && (_stream_conv2d_25_source_26_source_sel == 9);
  reg [_tmp_260-1:0] __tmp_261_1;
  assign _stream_conv2d_25_source_26_source_ram_rdata = (_stream_conv2d_25_source_26_source_sel == 9)? ram_w32_l4096_id7_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_336;
  assign stream_conv2d_25_source_26_data = __variable_wdata_336;
  reg [32-1:0] _stream_conv2d_25_source_26_source_pat_fsm_8;
  localparam _stream_conv2d_25_source_26_source_pat_fsm_8_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_26_source_pat_all_offset;
  assign _stream_conv2d_25_source_26_source_pat_all_offset = _stream_conv2d_25_source_26_source_offset_buf + _source_stream_conv2d_25_source_26_pat_cur_offset_0 + _source_stream_conv2d_25_source_26_pat_cur_offset_1 + _source_stream_conv2d_25_source_26_pat_cur_offset_2 + _source_stream_conv2d_25_source_26_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_25_source_27_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_27_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_27_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_27_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_27_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_27_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_27_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_27_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_27_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_27_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_27_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_27_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_27_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_27_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_27_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_27_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_27_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_27_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_27_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_27_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_27_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_27_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_27_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_27_pat_stride_buf_3;
  wire _set_flag_262;
  assign _set_flag_262 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l4096_id8_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_27_source_ram_renable && (_stream_conv2d_25_source_27_source_sel == 10))? _stream_conv2d_25_source_27_source_ram_raddr : 'hx;
  assign ram_w32_l4096_id8_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_27_source_ram_renable && (_stream_conv2d_25_source_27_source_sel == 10))? 1'd1 : 0;
  localparam _tmp_263 = 1;
  wire [_tmp_263-1:0] _tmp_264;
  assign _tmp_264 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_27_source_ram_renable && (_stream_conv2d_25_source_27_source_sel == 10);
  reg [_tmp_263-1:0] __tmp_264_1;
  assign _stream_conv2d_25_source_27_source_ram_rdata = (_stream_conv2d_25_source_27_source_sel == 10)? ram_w32_l4096_id8_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_337;
  assign stream_conv2d_25_source_27_data = __variable_wdata_337;
  reg [32-1:0] _stream_conv2d_25_source_27_source_pat_fsm_9;
  localparam _stream_conv2d_25_source_27_source_pat_fsm_9_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_27_source_pat_all_offset;
  assign _stream_conv2d_25_source_27_source_pat_all_offset = _stream_conv2d_25_source_27_source_offset_buf + _source_stream_conv2d_25_source_27_pat_cur_offset_0 + _source_stream_conv2d_25_source_27_pat_cur_offset_1 + _source_stream_conv2d_25_source_27_pat_cur_offset_2 + _source_stream_conv2d_25_source_27_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_25_source_28_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_28_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_28_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_28_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_28_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_28_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_28_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_28_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_28_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_28_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_28_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_28_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_28_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_28_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_28_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_28_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_28_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_28_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_28_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_28_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_28_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_28_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_28_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_28_pat_stride_buf_3;
  wire _set_flag_265;
  assign _set_flag_265 = conv2d_25_comp_fsm == 3;
  localparam _tmp_266 = 1;
  wire [_tmp_266-1:0] _tmp_267;
  assign _tmp_267 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_28_source_ram_renable && (_stream_conv2d_25_source_28_source_sel == 11);
  reg [_tmp_266-1:0] __tmp_267_1;
  assign _stream_conv2d_25_source_28_source_ram_rdata = (_stream_conv2d_25_source_28_source_sel == 11)? ram_w32_l8192_id0_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_338;
  assign stream_conv2d_25_source_28_data = __variable_wdata_338;
  reg [32-1:0] _stream_conv2d_25_source_28_source_pat_fsm_10;
  localparam _stream_conv2d_25_source_28_source_pat_fsm_10_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_28_source_pat_all_offset;
  assign _stream_conv2d_25_source_28_source_pat_all_offset = _stream_conv2d_25_source_28_source_offset_buf + _source_stream_conv2d_25_source_28_pat_cur_offset_0 + _source_stream_conv2d_25_source_28_pat_cur_offset_1 + _source_stream_conv2d_25_source_28_pat_cur_offset_2 + _source_stream_conv2d_25_source_28_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_25_source_29_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_29_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_29_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_29_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_29_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_29_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_29_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_29_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_29_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_29_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_29_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_29_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_29_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_29_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_29_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_29_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_29_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_29_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_29_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_29_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_29_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_29_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_29_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_29_pat_stride_buf_3;
  wire _set_flag_268;
  assign _set_flag_268 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l1024_id2_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_29_source_ram_renable && (_stream_conv2d_25_source_29_source_sel == 12))? _stream_conv2d_25_source_29_source_ram_raddr : 'hx;
  assign ram_w32_l1024_id2_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_29_source_ram_renable && (_stream_conv2d_25_source_29_source_sel == 12))? 1'd1 : 0;
  localparam _tmp_269 = 1;
  wire [_tmp_269-1:0] _tmp_270;
  assign _tmp_270 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_29_source_ram_renable && (_stream_conv2d_25_source_29_source_sel == 12);
  reg [_tmp_269-1:0] __tmp_270_1;
  assign _stream_conv2d_25_source_29_source_ram_rdata = (_stream_conv2d_25_source_29_source_sel == 12)? ram_w32_l1024_id2_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_564;
  assign stream_conv2d_25_source_29_data = __variable_wdata_564;
  reg [32-1:0] _stream_conv2d_25_source_29_source_pat_fsm_11;
  localparam _stream_conv2d_25_source_29_source_pat_fsm_11_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_29_source_pat_all_offset;
  assign _stream_conv2d_25_source_29_source_pat_all_offset = _stream_conv2d_25_source_29_source_offset_buf + _source_stream_conv2d_25_source_29_pat_cur_offset_0 + _source_stream_conv2d_25_source_29_pat_cur_offset_1 + _source_stream_conv2d_25_source_29_pat_cur_offset_2 + _source_stream_conv2d_25_source_29_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_25_source_30_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_30_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_30_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_30_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_30_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_30_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_30_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_30_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_30_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_30_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_30_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_30_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_30_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_30_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_30_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_30_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_30_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_30_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_30_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_30_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_30_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_30_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_30_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_30_pat_stride_buf_3;
  wire _set_flag_271;
  assign _set_flag_271 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l1024_id3_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_30_source_ram_renable && (_stream_conv2d_25_source_30_source_sel == 13))? _stream_conv2d_25_source_30_source_ram_raddr : 'hx;
  assign ram_w32_l1024_id3_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_30_source_ram_renable && (_stream_conv2d_25_source_30_source_sel == 13))? 1'd1 : 0;
  localparam _tmp_272 = 1;
  wire [_tmp_272-1:0] _tmp_273;
  assign _tmp_273 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_30_source_ram_renable && (_stream_conv2d_25_source_30_source_sel == 13);
  reg [_tmp_272-1:0] __tmp_273_1;
  assign _stream_conv2d_25_source_30_source_ram_rdata = (_stream_conv2d_25_source_30_source_sel == 13)? ram_w32_l1024_id3_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_565;
  assign stream_conv2d_25_source_30_data = __variable_wdata_565;
  reg [32-1:0] _stream_conv2d_25_source_30_source_pat_fsm_12;
  localparam _stream_conv2d_25_source_30_source_pat_fsm_12_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_30_source_pat_all_offset;
  assign _stream_conv2d_25_source_30_source_pat_all_offset = _stream_conv2d_25_source_30_source_offset_buf + _source_stream_conv2d_25_source_30_pat_cur_offset_0 + _source_stream_conv2d_25_source_30_pat_cur_offset_1 + _source_stream_conv2d_25_source_30_pat_cur_offset_2 + _source_stream_conv2d_25_source_30_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_25_source_31_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_31_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_31_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_31_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_31_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_31_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_31_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_31_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_31_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_31_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_31_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_31_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_31_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_31_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_31_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_31_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_31_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_31_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_31_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_31_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_31_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_31_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_31_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_31_pat_stride_buf_3;
  wire _set_flag_274;
  assign _set_flag_274 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l1024_id4_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_31_source_ram_renable && (_stream_conv2d_25_source_31_source_sel == 14))? _stream_conv2d_25_source_31_source_ram_raddr : 'hx;
  assign ram_w32_l1024_id4_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_31_source_ram_renable && (_stream_conv2d_25_source_31_source_sel == 14))? 1'd1 : 0;
  localparam _tmp_275 = 1;
  wire [_tmp_275-1:0] _tmp_276;
  assign _tmp_276 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_31_source_ram_renable && (_stream_conv2d_25_source_31_source_sel == 14);
  reg [_tmp_275-1:0] __tmp_276_1;
  assign _stream_conv2d_25_source_31_source_ram_rdata = (_stream_conv2d_25_source_31_source_sel == 14)? ram_w32_l1024_id4_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_566;
  assign stream_conv2d_25_source_31_data = __variable_wdata_566;
  reg [32-1:0] _stream_conv2d_25_source_31_source_pat_fsm_13;
  localparam _stream_conv2d_25_source_31_source_pat_fsm_13_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_31_source_pat_all_offset;
  assign _stream_conv2d_25_source_31_source_pat_all_offset = _stream_conv2d_25_source_31_source_offset_buf + _source_stream_conv2d_25_source_31_pat_cur_offset_0 + _source_stream_conv2d_25_source_31_pat_cur_offset_1 + _source_stream_conv2d_25_source_31_pat_cur_offset_2 + _source_stream_conv2d_25_source_31_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_25_source_32_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_32_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_32_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_32_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_32_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_32_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_32_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_32_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_32_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_32_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_32_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_32_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_32_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_32_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_32_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_32_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_32_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_32_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_32_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_32_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_32_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_32_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_32_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_32_pat_stride_buf_3;
  wire _set_flag_277;
  assign _set_flag_277 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l1024_id5_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_32_source_ram_renable && (_stream_conv2d_25_source_32_source_sel == 15))? _stream_conv2d_25_source_32_source_ram_raddr : 'hx;
  assign ram_w32_l1024_id5_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_32_source_ram_renable && (_stream_conv2d_25_source_32_source_sel == 15))? 1'd1 : 0;
  localparam _tmp_278 = 1;
  wire [_tmp_278-1:0] _tmp_279;
  assign _tmp_279 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_32_source_ram_renable && (_stream_conv2d_25_source_32_source_sel == 15);
  reg [_tmp_278-1:0] __tmp_279_1;
  assign _stream_conv2d_25_source_32_source_ram_rdata = (_stream_conv2d_25_source_32_source_sel == 15)? ram_w32_l1024_id5_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_567;
  assign stream_conv2d_25_source_32_data = __variable_wdata_567;
  reg [32-1:0] _stream_conv2d_25_source_32_source_pat_fsm_14;
  localparam _stream_conv2d_25_source_32_source_pat_fsm_14_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_32_source_pat_all_offset;
  assign _stream_conv2d_25_source_32_source_pat_all_offset = _stream_conv2d_25_source_32_source_offset_buf + _source_stream_conv2d_25_source_32_pat_cur_offset_0 + _source_stream_conv2d_25_source_32_pat_cur_offset_1 + _source_stream_conv2d_25_source_32_pat_cur_offset_2 + _source_stream_conv2d_25_source_32_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_25_source_33_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_33_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_33_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_33_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_33_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_33_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_33_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_33_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_33_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_33_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_33_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_33_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_33_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_33_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_33_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_33_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_33_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_33_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_33_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_33_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_33_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_33_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_33_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_33_pat_stride_buf_3;
  wire _set_flag_280;
  assign _set_flag_280 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l1024_id6_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_33_source_ram_renable && (_stream_conv2d_25_source_33_source_sel == 16))? _stream_conv2d_25_source_33_source_ram_raddr : 'hx;
  assign ram_w32_l1024_id6_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_33_source_ram_renable && (_stream_conv2d_25_source_33_source_sel == 16))? 1'd1 : 0;
  localparam _tmp_281 = 1;
  wire [_tmp_281-1:0] _tmp_282;
  assign _tmp_282 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_33_source_ram_renable && (_stream_conv2d_25_source_33_source_sel == 16);
  reg [_tmp_281-1:0] __tmp_282_1;
  assign _stream_conv2d_25_source_33_source_ram_rdata = (_stream_conv2d_25_source_33_source_sel == 16)? ram_w32_l1024_id6_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_568;
  assign stream_conv2d_25_source_33_data = __variable_wdata_568;
  reg [32-1:0] _stream_conv2d_25_source_33_source_pat_fsm_15;
  localparam _stream_conv2d_25_source_33_source_pat_fsm_15_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_33_source_pat_all_offset;
  assign _stream_conv2d_25_source_33_source_pat_all_offset = _stream_conv2d_25_source_33_source_offset_buf + _source_stream_conv2d_25_source_33_pat_cur_offset_0 + _source_stream_conv2d_25_source_33_pat_cur_offset_1 + _source_stream_conv2d_25_source_33_pat_cur_offset_2 + _source_stream_conv2d_25_source_33_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_25_source_34_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_34_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_34_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_34_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_34_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_34_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_34_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_34_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_34_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_34_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_34_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_34_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_34_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_34_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_34_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_34_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_34_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_34_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_34_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_34_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_34_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_34_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_34_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_34_pat_stride_buf_3;
  wire _set_flag_283;
  assign _set_flag_283 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l1024_id7_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_34_source_ram_renable && (_stream_conv2d_25_source_34_source_sel == 17))? _stream_conv2d_25_source_34_source_ram_raddr : 'hx;
  assign ram_w32_l1024_id7_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_34_source_ram_renable && (_stream_conv2d_25_source_34_source_sel == 17))? 1'd1 : 0;
  localparam _tmp_284 = 1;
  wire [_tmp_284-1:0] _tmp_285;
  assign _tmp_285 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_34_source_ram_renable && (_stream_conv2d_25_source_34_source_sel == 17);
  reg [_tmp_284-1:0] __tmp_285_1;
  assign _stream_conv2d_25_source_34_source_ram_rdata = (_stream_conv2d_25_source_34_source_sel == 17)? ram_w32_l1024_id7_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_569;
  assign stream_conv2d_25_source_34_data = __variable_wdata_569;
  reg [32-1:0] _stream_conv2d_25_source_34_source_pat_fsm_16;
  localparam _stream_conv2d_25_source_34_source_pat_fsm_16_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_34_source_pat_all_offset;
  assign _stream_conv2d_25_source_34_source_pat_all_offset = _stream_conv2d_25_source_34_source_offset_buf + _source_stream_conv2d_25_source_34_pat_cur_offset_0 + _source_stream_conv2d_25_source_34_pat_cur_offset_1 + _source_stream_conv2d_25_source_34_pat_cur_offset_2 + _source_stream_conv2d_25_source_34_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_25_source_35_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_35_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_35_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_35_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_35_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_35_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_35_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_35_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_35_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_35_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_35_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_35_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_35_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_35_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_35_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_35_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_35_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_35_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_35_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_35_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_35_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_35_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_35_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_35_pat_stride_buf_3;
  wire _set_flag_286;
  assign _set_flag_286 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l1024_id8_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_35_source_ram_renable && (_stream_conv2d_25_source_35_source_sel == 18))? _stream_conv2d_25_source_35_source_ram_raddr : 'hx;
  assign ram_w32_l1024_id8_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_35_source_ram_renable && (_stream_conv2d_25_source_35_source_sel == 18))? 1'd1 : 0;
  localparam _tmp_287 = 1;
  wire [_tmp_287-1:0] _tmp_288;
  assign _tmp_288 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_35_source_ram_renable && (_stream_conv2d_25_source_35_source_sel == 18);
  reg [_tmp_287-1:0] __tmp_288_1;
  assign _stream_conv2d_25_source_35_source_ram_rdata = (_stream_conv2d_25_source_35_source_sel == 18)? ram_w32_l1024_id8_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_570;
  assign stream_conv2d_25_source_35_data = __variable_wdata_570;
  reg [32-1:0] _stream_conv2d_25_source_35_source_pat_fsm_17;
  localparam _stream_conv2d_25_source_35_source_pat_fsm_17_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_35_source_pat_all_offset;
  assign _stream_conv2d_25_source_35_source_pat_all_offset = _stream_conv2d_25_source_35_source_offset_buf + _source_stream_conv2d_25_source_35_pat_cur_offset_0 + _source_stream_conv2d_25_source_35_pat_cur_offset_1 + _source_stream_conv2d_25_source_35_pat_cur_offset_2 + _source_stream_conv2d_25_source_35_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_25_source_36_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_36_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_36_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_36_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_36_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_36_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_36_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_36_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_36_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_36_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_36_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_36_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_36_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_36_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_36_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_36_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_36_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_36_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_36_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_36_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_36_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_36_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_36_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_36_pat_stride_buf_3;
  wire _set_flag_289;
  assign _set_flag_289 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l1024_id9_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_36_source_ram_renable && (_stream_conv2d_25_source_36_source_sel == 19))? _stream_conv2d_25_source_36_source_ram_raddr : 'hx;
  assign ram_w32_l1024_id9_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_36_source_ram_renable && (_stream_conv2d_25_source_36_source_sel == 19))? 1'd1 : 0;
  localparam _tmp_290 = 1;
  wire [_tmp_290-1:0] _tmp_291;
  assign _tmp_291 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_36_source_ram_renable && (_stream_conv2d_25_source_36_source_sel == 19);
  reg [_tmp_290-1:0] __tmp_291_1;
  assign _stream_conv2d_25_source_36_source_ram_rdata = (_stream_conv2d_25_source_36_source_sel == 19)? ram_w32_l1024_id9_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_571;
  assign stream_conv2d_25_source_36_data = __variable_wdata_571;
  reg [32-1:0] _stream_conv2d_25_source_36_source_pat_fsm_18;
  localparam _stream_conv2d_25_source_36_source_pat_fsm_18_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_36_source_pat_all_offset;
  assign _stream_conv2d_25_source_36_source_pat_all_offset = _stream_conv2d_25_source_36_source_offset_buf + _source_stream_conv2d_25_source_36_pat_cur_offset_0 + _source_stream_conv2d_25_source_36_pat_cur_offset_1 + _source_stream_conv2d_25_source_36_pat_cur_offset_2 + _source_stream_conv2d_25_source_36_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_25_source_37_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_25_source_37_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_25_source_37_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_25_source_37_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_25_source_37_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_25_source_37_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_25_source_37_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_25_source_37_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_25_source_37_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_25_source_37_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_25_source_37_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_25_source_37_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_25_source_37_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_25_source_37_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_25_source_37_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_25_source_37_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_25_source_37_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_25_source_37_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_25_source_37_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_25_source_37_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_25_source_37_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_25_source_37_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_25_source_37_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_25_source_37_pat_stride_buf_3;
  wire _set_flag_292;
  assign _set_flag_292 = conv2d_25_comp_fsm == 3;
  assign ram_w32_l1024_id10_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_37_source_ram_renable && (_stream_conv2d_25_source_37_source_sel == 20))? _stream_conv2d_25_source_37_source_ram_raddr : 'hx;
  assign ram_w32_l1024_id10_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_37_source_ram_renable && (_stream_conv2d_25_source_37_source_sel == 20))? 1'd1 : 0;
  localparam _tmp_293 = 1;
  wire [_tmp_293-1:0] _tmp_294;
  assign _tmp_294 = _stream_conv2d_25_stream_oready && _stream_conv2d_25_source_37_source_ram_renable && (_stream_conv2d_25_source_37_source_sel == 20);
  reg [_tmp_293-1:0] __tmp_294_1;
  assign _stream_conv2d_25_source_37_source_ram_rdata = (_stream_conv2d_25_source_37_source_sel == 20)? ram_w32_l1024_id10_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_572;
  assign stream_conv2d_25_source_37_data = __variable_wdata_572;
  reg [32-1:0] _stream_conv2d_25_source_37_source_pat_fsm_19;
  localparam _stream_conv2d_25_source_37_source_pat_fsm_19_init = 0;
  wire [32-1:0] _stream_conv2d_25_source_37_source_pat_all_offset;
  assign _stream_conv2d_25_source_37_source_pat_all_offset = _stream_conv2d_25_source_37_source_offset_buf + _source_stream_conv2d_25_source_37_pat_cur_offset_0 + _source_stream_conv2d_25_source_37_pat_cur_offset_1 + _source_stream_conv2d_25_source_37_pat_cur_offset_2 + _source_stream_conv2d_25_source_37_pat_cur_offset_3;
  wire _set_flag_295;
  assign _set_flag_295 = conv2d_25_comp_fsm == 3;
  reg _tmp_296;
  reg _tmp_297;
  reg _tmp_298;
  reg _tmp_299;
  reg _tmp_300;
  reg _tmp_301;
  reg _tmp_302;
  reg _tmp_303;
  reg _tmp_304;
  reg _tmp_305;
  reg _tmp_306;
  reg _tmp_307;
  reg _tmp_308;
  reg _tmp_309;
  reg _tmp_310;
  reg _tmp_311;
  reg _tmp_312;
  reg _tmp_313;
  reg _tmp_314;
  reg _tmp_315;
  reg _tmp_316;
  reg _tmp_317;
  reg _tmp_318;
  reg _tmp_319;
  reg _tmp_320;
  reg _tmp_321;
  reg _tmp_322;
  reg _tmp_323;
  reg _tmp_324;
  reg _tmp_325;
  reg _tmp_326;
  reg _tmp_327;
  reg _tmp_328;
  reg _tmp_329;
  reg _tmp_330;
  reg _tmp_331;
  localparam _tmp_332 = 33;
  wire [_tmp_332-1:0] _tmp_333;
  assign _tmp_333 = conv2d_25_stream_out_local + conv2d_25_out_page_comp_offset_buf;
  reg [_tmp_332-1:0] _tmp_334;
  reg [_tmp_332-1:0] _tmp_335;
  reg [_tmp_332-1:0] _tmp_336;
  reg [_tmp_332-1:0] _tmp_337;
  reg [_tmp_332-1:0] _tmp_338;
  reg [_tmp_332-1:0] _tmp_339;
  reg [_tmp_332-1:0] _tmp_340;
  reg [_tmp_332-1:0] _tmp_341;
  reg [_tmp_332-1:0] _tmp_342;
  reg [_tmp_332-1:0] _tmp_343;
  reg [_tmp_332-1:0] _tmp_344;
  reg [_tmp_332-1:0] _tmp_345;
  reg [_tmp_332-1:0] _tmp_346;
  reg [_tmp_332-1:0] _tmp_347;
  reg [_tmp_332-1:0] _tmp_348;
  reg [_tmp_332-1:0] _tmp_349;
  reg [_tmp_332-1:0] _tmp_350;
  reg [_tmp_332-1:0] _tmp_351;
  reg [_tmp_332-1:0] _tmp_352;
  reg [_tmp_332-1:0] _tmp_353;
  reg [_tmp_332-1:0] _tmp_354;
  reg [_tmp_332-1:0] _tmp_355;
  reg [_tmp_332-1:0] _tmp_356;
  reg [_tmp_332-1:0] _tmp_357;
  reg [_tmp_332-1:0] _tmp_358;
  reg [_tmp_332-1:0] _tmp_359;
  reg [_tmp_332-1:0] _tmp_360;
  reg [_tmp_332-1:0] _tmp_361;
  reg [_tmp_332-1:0] _tmp_362;
  reg [_tmp_332-1:0] _tmp_363;
  reg [_tmp_332-1:0] _tmp_364;
  reg [_tmp_332-1:0] _tmp_365;
  reg [_tmp_332-1:0] _tmp_366;
  reg [_tmp_332-1:0] _tmp_367;
  reg [_tmp_332-1:0] _tmp_368;
  reg [_tmp_332-1:0] _tmp_369;
  reg [32-1:0] _tmp_370;
  reg [32-1:0] _tmp_371;
  reg [32-1:0] _tmp_372;
  reg [32-1:0] _tmp_373;
  reg [32-1:0] _tmp_374;
  reg [32-1:0] _tmp_375;
  reg [32-1:0] _tmp_376;
  reg [32-1:0] _tmp_377;
  reg [32-1:0] _tmp_378;
  reg [32-1:0] _tmp_379;
  reg [32-1:0] _tmp_380;
  reg [32-1:0] _tmp_381;
  reg [32-1:0] _tmp_382;
  reg [32-1:0] _tmp_383;
  reg [32-1:0] _tmp_384;
  reg [32-1:0] _tmp_385;
  reg [32-1:0] _tmp_386;
  reg [32-1:0] _tmp_387;
  reg [32-1:0] _tmp_388;
  reg [32-1:0] _tmp_389;
  reg [32-1:0] _tmp_390;
  reg [32-1:0] _tmp_391;
  reg [32-1:0] _tmp_392;
  reg [32-1:0] _tmp_393;
  reg [32-1:0] _tmp_394;
  reg [32-1:0] _tmp_395;
  reg [32-1:0] _tmp_396;
  reg [32-1:0] _tmp_397;
  reg [32-1:0] _tmp_398;
  reg [32-1:0] _tmp_399;
  reg [32-1:0] _tmp_400;
  reg [32-1:0] _tmp_401;
  reg [32-1:0] _tmp_402;
  reg [32-1:0] _tmp_403;
  reg [32-1:0] _tmp_404;
  reg [32-1:0] _tmp_405;
  assign ram_w32_l1024_id1_0_addr = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_sink_50_sink_wenable && (_stream_conv2d_25_sink_50_sink_sel == 21))? _stream_conv2d_25_sink_50_sink_waddr : 'hx;
  assign ram_w32_l1024_id1_0_wdata = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_sink_50_sink_wenable && (_stream_conv2d_25_sink_50_sink_sel == 21))? _stream_conv2d_25_sink_50_sink_wdata : 'hx;
  assign ram_w32_l1024_id1_0_wenable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_sink_50_sink_wenable && (_stream_conv2d_25_sink_50_sink_sel == 21))? 1'd1 : 0;
  assign ram_w32_l1024_id1_0_enable = (_stream_conv2d_25_stream_oready && _stream_conv2d_25_sink_50_sink_wenable && (_stream_conv2d_25_sink_50_sink_sel == 21))? 1'd1 : 0;
  reg [32-1:0] _stream_conv2d_25_sink_50_sink_fsm_20;
  localparam _stream_conv2d_25_sink_50_sink_fsm_20_init = 0;
  wire _set_flag_406;
  assign _set_flag_406 = conv2d_25_comp_fsm == 4;
  assign _stream_conv2d_25_run_flag = (_set_flag_406)? 1 : 0;
  reg _tmp_407;
  reg _tmp_408;
  reg _tmp_409;
  assign _mul_4_source_stop = _mul_4_stream_oready && 1'd0;
  reg _tmp_410;
  reg _tmp_411;
  reg _tmp_412;
  reg _tmp_413;
  reg _tmp_414;
  reg _tmp_415;
  reg _tmp_416;
  reg _tmp_417;
  reg _tmp_418;
  reg _tmp_419;
  assign _mul_4_sink_start = _tmp_419;
  reg _tmp_420;
  reg _tmp_421;
  reg _tmp_422;
  reg _tmp_423;
  reg _tmp_424;
  reg _tmp_425;
  reg _tmp_426;
  reg _tmp_427;
  reg _tmp_428;
  reg _tmp_429;
  assign _mul_4_sink_stop = _tmp_429;
  reg _tmp_430;
  reg _tmp_431;
  reg _tmp_432;
  reg _tmp_433;
  reg _tmp_434;
  reg _tmp_435;
  reg _tmp_436;
  reg _tmp_437;
  reg _tmp_438;
  reg _tmp_439;
  assign _mul_4_sink_busy = _tmp_439;
  reg _tmp_440;
  assign _mul_4_busy = _mul_4_source_busy || _mul_4_sink_busy || _mul_4_busy_reg;
  reg _tmp_441;
  reg _tmp_442;
  reg _tmp_443;
  assign _mul_5_source_stop = _mul_5_stream_oready && 1'd0;
  reg _tmp_444;
  reg _tmp_445;
  reg _tmp_446;
  reg _tmp_447;
  reg _tmp_448;
  reg _tmp_449;
  reg _tmp_450;
  reg _tmp_451;
  reg _tmp_452;
  reg _tmp_453;
  assign _mul_5_sink_start = _tmp_453;
  reg _tmp_454;
  reg _tmp_455;
  reg _tmp_456;
  reg _tmp_457;
  reg _tmp_458;
  reg _tmp_459;
  reg _tmp_460;
  reg _tmp_461;
  reg _tmp_462;
  reg _tmp_463;
  assign _mul_5_sink_stop = _tmp_463;
  reg _tmp_464;
  reg _tmp_465;
  reg _tmp_466;
  reg _tmp_467;
  reg _tmp_468;
  reg _tmp_469;
  reg _tmp_470;
  reg _tmp_471;
  reg _tmp_472;
  reg _tmp_473;
  assign _mul_5_sink_busy = _tmp_473;
  reg _tmp_474;
  assign _mul_5_busy = _mul_5_source_busy || _mul_5_sink_busy || _mul_5_busy_reg;
  reg _tmp_475;
  reg _tmp_476;
  reg _tmp_477;
  assign _mul_6_source_stop = _mul_6_stream_oready && 1'd0;
  reg _tmp_478;
  reg _tmp_479;
  reg _tmp_480;
  reg _tmp_481;
  reg _tmp_482;
  reg _tmp_483;
  reg _tmp_484;
  reg _tmp_485;
  reg _tmp_486;
  reg _tmp_487;
  assign _mul_6_sink_start = _tmp_487;
  reg _tmp_488;
  reg _tmp_489;
  reg _tmp_490;
  reg _tmp_491;
  reg _tmp_492;
  reg _tmp_493;
  reg _tmp_494;
  reg _tmp_495;
  reg _tmp_496;
  reg _tmp_497;
  assign _mul_6_sink_stop = _tmp_497;
  reg _tmp_498;
  reg _tmp_499;
  reg _tmp_500;
  reg _tmp_501;
  reg _tmp_502;
  reg _tmp_503;
  reg _tmp_504;
  reg _tmp_505;
  reg _tmp_506;
  reg _tmp_507;
  assign _mul_6_sink_busy = _tmp_507;
  reg _tmp_508;
  assign _mul_6_busy = _mul_6_source_busy || _mul_6_sink_busy || _mul_6_busy_reg;
  reg _tmp_509;
  reg _tmp_510;
  reg _tmp_511;
  assign _mul_7_source_stop = _mul_7_stream_oready && 1'd0;
  reg _tmp_512;
  reg _tmp_513;
  reg _tmp_514;
  reg _tmp_515;
  reg _tmp_516;
  reg _tmp_517;
  reg _tmp_518;
  reg _tmp_519;
  reg _tmp_520;
  reg _tmp_521;
  assign _mul_7_sink_start = _tmp_521;
  reg _tmp_522;
  reg _tmp_523;
  reg _tmp_524;
  reg _tmp_525;
  reg _tmp_526;
  reg _tmp_527;
  reg _tmp_528;
  reg _tmp_529;
  reg _tmp_530;
  reg _tmp_531;
  assign _mul_7_sink_stop = _tmp_531;
  reg _tmp_532;
  reg _tmp_533;
  reg _tmp_534;
  reg _tmp_535;
  reg _tmp_536;
  reg _tmp_537;
  reg _tmp_538;
  reg _tmp_539;
  reg _tmp_540;
  reg _tmp_541;
  assign _mul_7_sink_busy = _tmp_541;
  reg _tmp_542;
  assign _mul_7_busy = _mul_7_source_busy || _mul_7_sink_busy || _mul_7_busy_reg;
  reg _tmp_543;
  reg _tmp_544;
  reg _tmp_545;
  assign _mul_8_source_stop = _mul_8_stream_oready && 1'd0;
  reg _tmp_546;
  reg _tmp_547;
  reg _tmp_548;
  reg _tmp_549;
  reg _tmp_550;
  reg _tmp_551;
  reg _tmp_552;
  reg _tmp_553;
  reg _tmp_554;
  reg _tmp_555;
  assign _mul_8_sink_start = _tmp_555;
  reg _tmp_556;
  reg _tmp_557;
  reg _tmp_558;
  reg _tmp_559;
  reg _tmp_560;
  reg _tmp_561;
  reg _tmp_562;
  reg _tmp_563;
  reg _tmp_564;
  reg _tmp_565;
  assign _mul_8_sink_stop = _tmp_565;
  reg _tmp_566;
  reg _tmp_567;
  reg _tmp_568;
  reg _tmp_569;
  reg _tmp_570;
  reg _tmp_571;
  reg _tmp_572;
  reg _tmp_573;
  reg _tmp_574;
  reg _tmp_575;
  assign _mul_8_sink_busy = _tmp_575;
  reg _tmp_576;
  assign _mul_8_busy = _mul_8_source_busy || _mul_8_sink_busy || _mul_8_busy_reg;
  reg _tmp_577;
  reg _tmp_578;
  reg _tmp_579;
  assign _mul_9_source_stop = _mul_9_stream_oready && 1'd0;
  reg _tmp_580;
  reg _tmp_581;
  reg _tmp_582;
  reg _tmp_583;
  reg _tmp_584;
  reg _tmp_585;
  reg _tmp_586;
  reg _tmp_587;
  reg _tmp_588;
  reg _tmp_589;
  assign _mul_9_sink_start = _tmp_589;
  reg _tmp_590;
  reg _tmp_591;
  reg _tmp_592;
  reg _tmp_593;
  reg _tmp_594;
  reg _tmp_595;
  reg _tmp_596;
  reg _tmp_597;
  reg _tmp_598;
  reg _tmp_599;
  assign _mul_9_sink_stop = _tmp_599;
  reg _tmp_600;
  reg _tmp_601;
  reg _tmp_602;
  reg _tmp_603;
  reg _tmp_604;
  reg _tmp_605;
  reg _tmp_606;
  reg _tmp_607;
  reg _tmp_608;
  reg _tmp_609;
  assign _mul_9_sink_busy = _tmp_609;
  reg _tmp_610;
  assign _mul_9_busy = _mul_9_source_busy || _mul_9_sink_busy || _mul_9_busy_reg;
  reg _tmp_611;
  reg _tmp_612;
  reg _tmp_613;
  assign _mul_10_source_stop = _mul_10_stream_oready && 1'd0;
  reg _tmp_614;
  reg _tmp_615;
  reg _tmp_616;
  reg _tmp_617;
  reg _tmp_618;
  reg _tmp_619;
  reg _tmp_620;
  reg _tmp_621;
  reg _tmp_622;
  reg _tmp_623;
  assign _mul_10_sink_start = _tmp_623;
  reg _tmp_624;
  reg _tmp_625;
  reg _tmp_626;
  reg _tmp_627;
  reg _tmp_628;
  reg _tmp_629;
  reg _tmp_630;
  reg _tmp_631;
  reg _tmp_632;
  reg _tmp_633;
  assign _mul_10_sink_stop = _tmp_633;
  reg _tmp_634;
  reg _tmp_635;
  reg _tmp_636;
  reg _tmp_637;
  reg _tmp_638;
  reg _tmp_639;
  reg _tmp_640;
  reg _tmp_641;
  reg _tmp_642;
  reg _tmp_643;
  assign _mul_10_sink_busy = _tmp_643;
  reg _tmp_644;
  assign _mul_10_busy = _mul_10_source_busy || _mul_10_sink_busy || _mul_10_busy_reg;
  reg _tmp_645;
  reg _tmp_646;
  reg _tmp_647;
  assign _mul_11_source_stop = _mul_11_stream_oready && 1'd0;
  reg _tmp_648;
  reg _tmp_649;
  reg _tmp_650;
  reg _tmp_651;
  reg _tmp_652;
  reg _tmp_653;
  reg _tmp_654;
  reg _tmp_655;
  reg _tmp_656;
  reg _tmp_657;
  assign _mul_11_sink_start = _tmp_657;
  reg _tmp_658;
  reg _tmp_659;
  reg _tmp_660;
  reg _tmp_661;
  reg _tmp_662;
  reg _tmp_663;
  reg _tmp_664;
  reg _tmp_665;
  reg _tmp_666;
  reg _tmp_667;
  assign _mul_11_sink_stop = _tmp_667;
  reg _tmp_668;
  reg _tmp_669;
  reg _tmp_670;
  reg _tmp_671;
  reg _tmp_672;
  reg _tmp_673;
  reg _tmp_674;
  reg _tmp_675;
  reg _tmp_676;
  reg _tmp_677;
  assign _mul_11_sink_busy = _tmp_677;
  reg _tmp_678;
  assign _mul_11_busy = _mul_11_source_busy || _mul_11_sink_busy || _mul_11_busy_reg;
  reg _tmp_679;
  reg _tmp_680;
  reg _tmp_681;
  assign _mul_12_source_stop = _mul_12_stream_oready && 1'd0;
  reg _tmp_682;
  reg _tmp_683;
  reg _tmp_684;
  reg _tmp_685;
  reg _tmp_686;
  reg _tmp_687;
  reg _tmp_688;
  reg _tmp_689;
  reg _tmp_690;
  reg _tmp_691;
  assign _mul_12_sink_start = _tmp_691;
  reg _tmp_692;
  reg _tmp_693;
  reg _tmp_694;
  reg _tmp_695;
  reg _tmp_696;
  reg _tmp_697;
  reg _tmp_698;
  reg _tmp_699;
  reg _tmp_700;
  reg _tmp_701;
  assign _mul_12_sink_stop = _tmp_701;
  reg _tmp_702;
  reg _tmp_703;
  reg _tmp_704;
  reg _tmp_705;
  reg _tmp_706;
  reg _tmp_707;
  reg _tmp_708;
  reg _tmp_709;
  reg _tmp_710;
  reg _tmp_711;
  assign _mul_12_sink_busy = _tmp_711;
  reg _tmp_712;
  assign _mul_12_busy = _mul_12_source_busy || _mul_12_sink_busy || _mul_12_busy_reg;
  reg _tmp_713;
  reg _tmp_714;
  reg _tmp_715;
  assign _add_tree_2_source_stop = _add_tree_2_stream_oready && 1'd0;
  reg _tmp_716;
  reg _tmp_717;
  reg _tmp_718;
  reg _tmp_719;
  assign _add_tree_2_sink_start = _tmp_719;
  reg _tmp_720;
  reg _tmp_721;
  reg _tmp_722;
  reg _tmp_723;
  assign _add_tree_2_sink_stop = _tmp_723;
  reg _tmp_724;
  reg _tmp_725;
  reg _tmp_726;
  reg _tmp_727;
  assign _add_tree_2_sink_busy = _tmp_727;
  reg _tmp_728;
  assign _add_tree_2_busy = _add_tree_2_source_busy || _add_tree_2_sink_busy || _add_tree_2_busy_reg;
  reg _tmp_729;
  reg _tmp_730;
  reg _tmp_731;
  reg _tmp_732;
  reg _tmp_733;
  reg _tmp_734;
  reg _tmp_735;
  reg _tmp_736;
  reg _tmp_737;
  reg _tmp_738;
  assign _acc_1_source_stop = _acc_1_stream_oready && 1'd0;
  reg _tmp_739;
  reg _tmp_740;
  reg _tmp_741;
  reg _tmp_742;
  reg _tmp_743;
  reg _tmp_744;
  reg _tmp_745;
  assign _acc_1_sink_start = _tmp_745;
  reg _tmp_746;
  reg _tmp_747;
  reg _tmp_748;
  reg _tmp_749;
  reg _tmp_750;
  reg _tmp_751;
  reg _tmp_752;
  assign _acc_1_sink_stop = _tmp_752;
  reg _tmp_753;
  reg _tmp_754;
  reg _tmp_755;
  reg _tmp_756;
  reg _tmp_757;
  reg _tmp_758;
  reg _tmp_759;
  assign _acc_1_sink_busy = _tmp_759;
  reg _tmp_760;
  assign _acc_1_busy = _acc_1_source_busy || _acc_1_sink_busy || _acc_1_busy_reg;
  reg _tmp_761;
  reg _tmp_762;
  reg _tmp_763;
  assign _mul_rshift_round_clip_3_source_stop = _mul_rshift_round_clip_3_stream_oready && 1'd0;
  reg _tmp_764;
  reg _tmp_765;
  reg _tmp_766;
  reg _tmp_767;
  reg _tmp_768;
  reg _tmp_769;
  reg _tmp_770;
  reg _tmp_771;
  reg _tmp_772;
  reg _tmp_773;
  assign _mul_rshift_round_clip_3_sink_start = _tmp_773;
  reg _tmp_774;
  reg _tmp_775;
  reg _tmp_776;
  reg _tmp_777;
  reg _tmp_778;
  reg _tmp_779;
  reg _tmp_780;
  reg _tmp_781;
  reg _tmp_782;
  reg _tmp_783;
  assign _mul_rshift_round_clip_3_sink_stop = _tmp_783;
  reg _tmp_784;
  reg _tmp_785;
  reg _tmp_786;
  reg _tmp_787;
  reg _tmp_788;
  reg _tmp_789;
  reg _tmp_790;
  reg _tmp_791;
  reg _tmp_792;
  reg _tmp_793;
  assign _mul_rshift_round_clip_3_sink_busy = _tmp_793;
  reg _tmp_794;
  assign _mul_rshift_round_clip_3_busy = _mul_rshift_round_clip_3_source_busy || _mul_rshift_round_clip_3_sink_busy || _mul_rshift_round_clip_3_busy_reg;
  reg _tmp_795;
  reg _tmp_796;
  reg _tmp_797;
  reg _tmp_798;
  reg _tmp_799;
  reg _tmp_800;
  reg [1-1:0] __variable_wdata_281;
  assign stream_conv2d_25__reduce_reset_data = __variable_wdata_281;
  reg _tmp_801;
  reg _tmp_802;
  reg _tmp_803;
  reg _tmp_804;
  assign _stream_conv2d_25_source_stop = _stream_conv2d_25_stream_oready && (_stream_conv2d_25_source_11_idle && _stream_conv2d_25_source_13_idle && _stream_conv2d_25_source_15_idle && _stream_conv2d_25_source_20_idle && _stream_conv2d_25_source_21_idle && _stream_conv2d_25_source_22_idle && _stream_conv2d_25_source_23_idle && _stream_conv2d_25_source_24_idle && _stream_conv2d_25_source_25_idle && _stream_conv2d_25_source_26_idle && _stream_conv2d_25_source_27_idle && _stream_conv2d_25_source_28_idle && _stream_conv2d_25_source_29_idle && _stream_conv2d_25_source_30_idle && _stream_conv2d_25_source_31_idle && _stream_conv2d_25_source_32_idle && _stream_conv2d_25_source_33_idle && _stream_conv2d_25_source_34_idle && _stream_conv2d_25_source_35_idle && _stream_conv2d_25_source_36_idle && _stream_conv2d_25_source_37_idle && _stream_conv2d_25_source_7_idle && _stream_conv2d_25_source_9_idle && (_stream_conv2d_25_fsm == 3));
  localparam _tmp_805 = 1;
  wire [_tmp_805-1:0] _tmp_806;
  assign _tmp_806 = _stream_conv2d_25_source_11_idle && _stream_conv2d_25_source_13_idle && _stream_conv2d_25_source_15_idle && _stream_conv2d_25_source_20_idle && _stream_conv2d_25_source_21_idle && _stream_conv2d_25_source_22_idle && _stream_conv2d_25_source_23_idle && _stream_conv2d_25_source_24_idle && _stream_conv2d_25_source_25_idle && _stream_conv2d_25_source_26_idle && _stream_conv2d_25_source_27_idle && _stream_conv2d_25_source_28_idle && _stream_conv2d_25_source_29_idle && _stream_conv2d_25_source_30_idle && _stream_conv2d_25_source_31_idle && _stream_conv2d_25_source_32_idle && _stream_conv2d_25_source_33_idle && _stream_conv2d_25_source_34_idle && _stream_conv2d_25_source_35_idle && _stream_conv2d_25_source_36_idle && _stream_conv2d_25_source_37_idle && _stream_conv2d_25_source_7_idle && _stream_conv2d_25_source_9_idle && (_stream_conv2d_25_fsm == 3);
  reg [_tmp_805-1:0] _tmp_807;
  localparam _tmp_808 = 1;
  wire [_tmp_808-1:0] _tmp_809;
  assign _tmp_809 = _stream_conv2d_25_source_11_idle && _stream_conv2d_25_source_13_idle && _stream_conv2d_25_source_15_idle && _stream_conv2d_25_source_20_idle && _stream_conv2d_25_source_21_idle && _stream_conv2d_25_source_22_idle && _stream_conv2d_25_source_23_idle && _stream_conv2d_25_source_24_idle && _stream_conv2d_25_source_25_idle && _stream_conv2d_25_source_26_idle && _stream_conv2d_25_source_27_idle && _stream_conv2d_25_source_28_idle && _stream_conv2d_25_source_29_idle && _stream_conv2d_25_source_30_idle && _stream_conv2d_25_source_31_idle && _stream_conv2d_25_source_32_idle && _stream_conv2d_25_source_33_idle && _stream_conv2d_25_source_34_idle && _stream_conv2d_25_source_35_idle && _stream_conv2d_25_source_36_idle && _stream_conv2d_25_source_37_idle && _stream_conv2d_25_source_7_idle && _stream_conv2d_25_source_9_idle && (_stream_conv2d_25_fsm == 3);
  reg [_tmp_808-1:0] _tmp_810;
  reg _tmp_811;
  reg _tmp_812;
  reg _tmp_813;
  reg _tmp_814;
  reg _tmp_815;
  reg _tmp_816;
  reg _tmp_817;
  reg _tmp_818;
  reg _tmp_819;
  reg _tmp_820;
  reg _tmp_821;
  reg _tmp_822;
  reg _tmp_823;
  reg _tmp_824;
  reg _tmp_825;
  reg _tmp_826;
  reg _tmp_827;
  reg _tmp_828;
  reg _tmp_829;
  reg _tmp_830;
  reg _tmp_831;
  reg _tmp_832;
  reg _tmp_833;
  reg _tmp_834;
  reg _tmp_835;
  reg _tmp_836;
  reg _tmp_837;
  reg _tmp_838;
  reg _tmp_839;
  reg _tmp_840;
  reg _tmp_841;
  reg _tmp_842;
  reg _tmp_843;
  reg _tmp_844;
  reg _tmp_845;
  reg _tmp_846;
  assign _stream_conv2d_25_sink_start = _tmp_846;
  reg _tmp_847;
  reg _tmp_848;
  reg _tmp_849;
  reg _tmp_850;
  reg _tmp_851;
  reg _tmp_852;
  reg _tmp_853;
  reg _tmp_854;
  reg _tmp_855;
  reg _tmp_856;
  reg _tmp_857;
  reg _tmp_858;
  reg _tmp_859;
  reg _tmp_860;
  reg _tmp_861;
  reg _tmp_862;
  reg _tmp_863;
  reg _tmp_864;
  reg _tmp_865;
  reg _tmp_866;
  reg _tmp_867;
  reg _tmp_868;
  reg _tmp_869;
  reg _tmp_870;
  reg _tmp_871;
  reg _tmp_872;
  reg _tmp_873;
  reg _tmp_874;
  reg _tmp_875;
  reg _tmp_876;
  reg _tmp_877;
  reg _tmp_878;
  reg _tmp_879;
  reg _tmp_880;
  reg _tmp_881;
  reg _tmp_882;
  assign _stream_conv2d_25_sink_stop = _tmp_882;
  reg _tmp_883;
  reg _tmp_884;
  reg _tmp_885;
  reg _tmp_886;
  reg _tmp_887;
  reg _tmp_888;
  reg _tmp_889;
  reg _tmp_890;
  reg _tmp_891;
  reg _tmp_892;
  reg _tmp_893;
  reg _tmp_894;
  reg _tmp_895;
  reg _tmp_896;
  reg _tmp_897;
  reg _tmp_898;
  reg _tmp_899;
  reg _tmp_900;
  reg _tmp_901;
  reg _tmp_902;
  reg _tmp_903;
  reg _tmp_904;
  reg _tmp_905;
  reg _tmp_906;
  reg _tmp_907;
  reg _tmp_908;
  reg _tmp_909;
  reg _tmp_910;
  reg _tmp_911;
  reg _tmp_912;
  reg _tmp_913;
  reg _tmp_914;
  reg _tmp_915;
  reg _tmp_916;
  reg _tmp_917;
  reg _tmp_918;
  assign _stream_conv2d_25_sink_busy = _tmp_918;
  reg _tmp_919;
  assign _stream_conv2d_25_busy = _stream_conv2d_25_source_busy || _stream_conv2d_25_sink_busy || _stream_conv2d_25_busy_reg;
  wire conv2d_25_dma_out_mask_0;
  assign conv2d_25_dma_out_mask_0 = conv2d_25_out_row_count + 0 >= cparam_conv2d_25_out_num_row;
  wire [32-1:0] mask_addr_shifted_920;
  assign mask_addr_shifted_920 = conv2d_25_objaddr + (conv2d_25_out_base_offset + cparam_conv2d_25_out_offset_values_0) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_921;
  assign mask_addr_masked_921 = mask_addr_shifted_920 << 2;
  reg [32-1:0] _maxi_write_req_fsm;
  localparam _maxi_write_req_fsm_init = 0;
  reg [33-1:0] _maxi_write_cur_global_size;
  reg _maxi_write_cont;
  wire [8-1:0] pack_write_req_op_sel_922;
  wire [32-1:0] pack_write_req_local_addr_923;
  wire [32-1:0] pack_write_req_local_stride_924;
  wire [33-1:0] pack_write_req_size_925;
  wire [32-1:0] pack_write_req_local_blocksize_926;
  assign pack_write_req_op_sel_922 = _maxi_write_op_sel;
  assign pack_write_req_local_addr_923 = _maxi_write_local_addr;
  assign pack_write_req_local_stride_924 = _maxi_write_local_stride;
  assign pack_write_req_size_925 = _maxi_write_local_size;
  assign pack_write_req_local_blocksize_926 = _maxi_write_local_blocksize;
  wire [137-1:0] pack_write_req_packed_927;
  assign pack_write_req_packed_927 = { pack_write_req_op_sel_922, pack_write_req_local_addr_923, pack_write_req_local_stride_924, pack_write_req_size_925, pack_write_req_local_blocksize_926 };
  localparam _tmp_928 = 1;
  wire [_tmp_928-1:0] _tmp_929;
  assign _tmp_929 = !_maxi_write_req_fifo_almost_full;
  reg [_tmp_928-1:0] __tmp_929_1;
  wire [32-1:0] mask_addr_shifted_930;
  assign mask_addr_shifted_930 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_931;
  assign mask_addr_masked_931 = mask_addr_shifted_930 << 2;
  wire [32-1:0] mask_addr_shifted_932;
  assign mask_addr_shifted_932 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_933;
  assign mask_addr_masked_933 = mask_addr_shifted_932 << 2;
  wire [32-1:0] mask_addr_shifted_934;
  assign mask_addr_shifted_934 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_935;
  assign mask_addr_masked_935 = mask_addr_shifted_934 << 2;
  wire [32-1:0] mask_addr_shifted_936;
  assign mask_addr_shifted_936 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_937;
  assign mask_addr_masked_937 = mask_addr_shifted_936 << 2;
  wire [32-1:0] mask_addr_shifted_938;
  assign mask_addr_shifted_938 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_939;
  assign mask_addr_masked_939 = mask_addr_shifted_938 << 2;
  wire [32-1:0] mask_addr_shifted_940;
  assign mask_addr_shifted_940 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_941;
  assign mask_addr_masked_941 = mask_addr_shifted_940 << 2;
  wire [8-1:0] pack_write_req_op_sel_942;
  wire [32-1:0] pack_write_req_local_addr_943;
  wire [32-1:0] pack_write_req_local_stride_944;
  wire [33-1:0] pack_write_req_size_945;
  wire [32-1:0] pack_write_req_local_blocksize_946;
  assign pack_write_req_op_sel_942 = _maxi_write_op_sel;
  assign pack_write_req_local_addr_943 = _maxi_write_local_addr;
  assign pack_write_req_local_stride_944 = _maxi_write_local_stride;
  assign pack_write_req_size_945 = _maxi_write_cur_global_size;
  assign pack_write_req_local_blocksize_946 = _maxi_write_local_blocksize;
  wire [137-1:0] pack_write_req_packed_947;
  assign pack_write_req_packed_947 = { pack_write_req_op_sel_942, pack_write_req_local_addr_943, pack_write_req_local_stride_944, pack_write_req_size_945, pack_write_req_local_blocksize_946 };
  assign _maxi_write_req_fifo_wdata = ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6))? pack_write_req_packed_947 : 
                                      ((_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full)? pack_write_req_packed_927 : 'hx;
  assign _maxi_write_req_fifo_enq = ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6))? (_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6) && !_maxi_write_req_fifo_almost_full : 
                                    ((_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full)? (_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full && !_maxi_write_req_fifo_almost_full : 0;
  localparam _tmp_948 = 1;
  wire [_tmp_948-1:0] _tmp_949;
  assign _tmp_949 = !_maxi_write_req_fifo_almost_full;
  reg [_tmp_948-1:0] __tmp_949_1;
  reg _maxi_waddr_cond_0_1;
  reg [32-1:0] _maxi_write_data_fsm;
  localparam _maxi_write_data_fsm_init = 0;
  reg [32-1:0] read_burst_fsm_24;
  localparam read_burst_fsm_24_init = 0;
  reg [10-1:0] read_burst_addr_950;
  reg [10-1:0] read_burst_stride_951;
  reg [33-1:0] read_burst_length_952;
  reg read_burst_rvalid_953;
  reg read_burst_rlast_954;
  assign ram_w32_l1024_id1_1_addr = ((read_burst_fsm_24 == 1) && (!read_burst_rvalid_953 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_addr_950 : 'hx;
  assign ram_w32_l1024_id1_1_enable = ((read_burst_fsm_24 == 1) && (!read_burst_rvalid_953 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 0;
  localparam _tmp_955 = 1;
  wire [_tmp_955-1:0] _tmp_956;
  assign _tmp_956 = (read_burst_fsm_24 == 1) && (!read_burst_rvalid_953 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_955-1:0] __tmp_956_1;
  wire [32-1:0] read_burst_rdata_957;
  assign read_burst_rdata_957 = ram_w32_l1024_id1_1_rdata;
  reg _maxi_wdata_cond_0_1;
  wire conv2d_25_update_filter;
  assign conv2d_25_update_filter = (cparam_conv2d_25_data_stationary == 0) && (conv2d_25_row_count >= cparam_conv2d_25_max_row_count) && (conv2d_25_bat_count >= cparam_conv2d_25_max_bat_count) || (cparam_conv2d_25_data_stationary == 1) && !cparam_conv2d_25_keep_filter;
  wire conv2d_25_update_act;
  assign conv2d_25_update_act = (cparam_conv2d_25_data_stationary == 1) && (conv2d_25_och_count >= cparam_conv2d_25_max_och_count) || (cparam_conv2d_25_data_stationary == 0);
  wire conv2d_25_mux_next_dma_flag_0;
  assign conv2d_25_mux_next_dma_flag_0 = (conv2d_25_row_select == 0)? (conv2d_25_row_count >= cparam_conv2d_25_max_row_count)? 1 : cparam_conv2d_25_dma_flag_conds_0 : 
                                         (conv2d_25_row_select == 1)? (conv2d_25_row_count >= cparam_conv2d_25_max_row_count)? 1 : cparam_conv2d_25_dma_flag_conds_2 : 
                                         (conv2d_25_row_select == 2)? (conv2d_25_row_count >= cparam_conv2d_25_max_row_count)? 1 : cparam_conv2d_25_dma_flag_conds_1 : 1'd0;
  wire conv2d_25_mux_next_dma_flag_1;
  assign conv2d_25_mux_next_dma_flag_1 = (conv2d_25_row_select == 0)? (conv2d_25_row_count >= cparam_conv2d_25_max_row_count)? 1 : cparam_conv2d_25_dma_flag_conds_1 : 
                                         (conv2d_25_row_select == 1)? (conv2d_25_row_count >= cparam_conv2d_25_max_row_count)? 1 : cparam_conv2d_25_dma_flag_conds_0 : 
                                         (conv2d_25_row_select == 2)? (conv2d_25_row_count >= cparam_conv2d_25_max_row_count)? 1 : cparam_conv2d_25_dma_flag_conds_2 : 1'd0;
  wire conv2d_25_mux_next_dma_flag_2;
  assign conv2d_25_mux_next_dma_flag_2 = (conv2d_25_row_select == 0)? (conv2d_25_row_count >= cparam_conv2d_25_max_row_count)? 1 : cparam_conv2d_25_dma_flag_conds_2 : 
                                         (conv2d_25_row_select == 1)? (conv2d_25_row_count >= cparam_conv2d_25_max_row_count)? 1 : cparam_conv2d_25_dma_flag_conds_1 : 
                                         (conv2d_25_row_select == 2)? (conv2d_25_row_count >= cparam_conv2d_25_max_row_count)? 1 : cparam_conv2d_25_dma_flag_conds_0 : 1'd0;
  reg [32-1:0] max_pool_serial_27_objaddr;
  reg [32-1:0] max_pool_serial_27_arg_objaddr_0;
  reg [32-1:0] control_max_pool_serial_27;
  localparam control_max_pool_serial_27_init = 0;
  reg _control_max_pool_serial_27_called;
  wire signed [32-1:0] max_pool_serial_27_act_base_offset;
  reg signed [32-1:0] max_pool_serial_27_act_base_offset_row;
  reg signed [32-1:0] max_pool_serial_27_act_base_offset_bat;
  assign max_pool_serial_27_act_base_offset = max_pool_serial_27_act_base_offset_row + max_pool_serial_27_act_base_offset_bat;
  wire signed [32-1:0] max_pool_serial_27_out_base_offset;
  reg signed [32-1:0] max_pool_serial_27_out_base_offset_row;
  reg signed [32-1:0] max_pool_serial_27_out_base_offset_bat;
  assign max_pool_serial_27_out_base_offset = max_pool_serial_27_out_base_offset_row + max_pool_serial_27_out_base_offset_bat;
  reg [32-1:0] max_pool_serial_27_col_count;
  reg [32-1:0] max_pool_serial_27_row_count;
  reg [32-1:0] max_pool_serial_27_bat_count;
  reg [32-1:0] max_pool_serial_27_prev_row_count;
  reg [32-1:0] max_pool_serial_27_prev_bat_count;
  reg [32-1:0] max_pool_serial_27_stream_act_local;
  reg [32-1:0] max_pool_serial_27_stream_out_local;
  reg max_pool_serial_27_act_page;
  reg [32-1:0] max_pool_serial_27_act_page_comp_offset;
  reg [32-1:0] max_pool_serial_27_act_page_dma_offset;
  reg max_pool_serial_27_out_page;
  reg [32-1:0] max_pool_serial_27_out_page_comp_offset;
  reg [32-1:0] max_pool_serial_27_out_page_dma_offset;
  reg max_pool_serial_27_skip_read_act;
  reg max_pool_serial_27_skip_comp;
  reg max_pool_serial_27_skip_write_out;
  reg [32-1:0] max_pool_serial_27_comp_count;
  reg [32-1:0] max_pool_serial_27_out_count;
  wire max_pool_serial_27_dma_pad_mask_0;
  assign max_pool_serial_27_dma_pad_mask_0 = (max_pool_serial_27_row_count + 0 < cparam_max_pool_serial_27_pad_row_top) || (max_pool_serial_27_row_count + 0 >= cparam_max_pool_serial_27_act_num_row + cparam_max_pool_serial_27_pad_row_top);
  wire max_pool_serial_27_dma_pad_mask_1;
  assign max_pool_serial_27_dma_pad_mask_1 = (max_pool_serial_27_row_count + 1 < cparam_max_pool_serial_27_pad_row_top) || (max_pool_serial_27_row_count + 1 >= cparam_max_pool_serial_27_act_num_row + cparam_max_pool_serial_27_pad_row_top);
  wire [32-1:0] mask_addr_shifted_958;
  assign mask_addr_shifted_958 = max_pool_serial_27_arg_objaddr_0 + (max_pool_serial_27_act_base_offset + cparam_max_pool_serial_27_act_offset_values_0) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_959;
  assign mask_addr_masked_959 = mask_addr_shifted_958 << 2;
  reg [32-1:0] write_burst_fsm_25;
  localparam write_burst_fsm_25_init = 0;
  reg [15-1:0] write_burst_addr_960;
  reg [15-1:0] write_burst_stride_961;
  reg [33-1:0] write_burst_length_962;
  reg write_burst_done_963;
  assign ram_w32_l32768_id0_1_addr = ((write_burst_fsm_25 == 1) && _maxi_rvalid_sb_0)? write_burst_addr_960 : 'hx;
  assign ram_w32_l32768_id0_1_wdata = ((write_burst_fsm_25 == 1) && _maxi_rvalid_sb_0)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l32768_id0_1_wenable = ((write_burst_fsm_25 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w32_l32768_id0_1_enable = ((write_burst_fsm_25 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [32-1:0] mask_addr_shifted_964;
  assign mask_addr_shifted_964 = max_pool_serial_27_arg_objaddr_0 + (max_pool_serial_27_act_base_offset + cparam_max_pool_serial_27_act_offset_values_1) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_965;
  assign mask_addr_masked_965 = mask_addr_shifted_964 << 2;
  reg [32-1:0] max_pool_serial_27_comp_fsm;
  localparam max_pool_serial_27_comp_fsm_init = 0;
  reg [32-1:0] max_pool_serial_27_act_page_comp_offset_buf;
  reg [32-1:0] max_pool_serial_27_out_page_comp_offset_buf;
  reg [32-1:0] max_pool_serial_27_row_count_buf;
  wire max_pool_serial_27_stream_pad_mask_0_0;
  assign max_pool_serial_27_stream_pad_mask_0_0 = (max_pool_serial_27_col_count + 0 < cparam_max_pool_serial_27_pad_col_left) || (max_pool_serial_27_col_count + 0 >= cparam_max_pool_serial_27_act_num_col + cparam_max_pool_serial_27_pad_col_left) || (max_pool_serial_27_row_count_buf + 0 < cparam_max_pool_serial_27_pad_row_top) || (max_pool_serial_27_row_count_buf + 0 >= cparam_max_pool_serial_27_act_num_row + cparam_max_pool_serial_27_pad_row_top);
  wire max_pool_serial_27_stream_pad_mask_0_1;
  assign max_pool_serial_27_stream_pad_mask_0_1 = (max_pool_serial_27_col_count + 1 < cparam_max_pool_serial_27_pad_col_left) || (max_pool_serial_27_col_count + 1 >= cparam_max_pool_serial_27_act_num_col + cparam_max_pool_serial_27_pad_col_left) || (max_pool_serial_27_row_count_buf + 0 < cparam_max_pool_serial_27_pad_row_top) || (max_pool_serial_27_row_count_buf + 0 >= cparam_max_pool_serial_27_act_num_row + cparam_max_pool_serial_27_pad_row_top);
  wire max_pool_serial_27_stream_pad_mask_1_0;
  assign max_pool_serial_27_stream_pad_mask_1_0 = (max_pool_serial_27_col_count + 0 < cparam_max_pool_serial_27_pad_col_left) || (max_pool_serial_27_col_count + 0 >= cparam_max_pool_serial_27_act_num_col + cparam_max_pool_serial_27_pad_col_left) || (max_pool_serial_27_row_count_buf + 1 < cparam_max_pool_serial_27_pad_row_top) || (max_pool_serial_27_row_count_buf + 1 >= cparam_max_pool_serial_27_act_num_row + cparam_max_pool_serial_27_pad_row_top);
  wire max_pool_serial_27_stream_pad_mask_1_1;
  assign max_pool_serial_27_stream_pad_mask_1_1 = (max_pool_serial_27_col_count + 1 < cparam_max_pool_serial_27_pad_col_left) || (max_pool_serial_27_col_count + 1 >= cparam_max_pool_serial_27_act_num_col + cparam_max_pool_serial_27_pad_col_left) || (max_pool_serial_27_row_count_buf + 1 < cparam_max_pool_serial_27_pad_row_top) || (max_pool_serial_27_row_count_buf + 1 >= cparam_max_pool_serial_27_act_num_row + cparam_max_pool_serial_27_pad_row_top);
  reg [4-1:0] max_pool_serial_27_stream_pad_masks;
  wire [3-1:0] stream_max_pool_serial_27_parameter_0_data;
  wire [32-1:0] stream_max_pool_serial_27_source_1_data;
  wire [4-1:0] stream_max_pool_serial_27_parameter_2_data;
  wire [1-1:0] stream_max_pool_serial_27__reduce_reset_data;
  reg __stream_max_pool_serial_27_stream_ivalid_1;
  reg __stream_max_pool_serial_27_stream_ivalid_2;
  reg __stream_max_pool_serial_27_stream_ivalid_3;
  reg __stream_max_pool_serial_27_stream_ivalid_4;
  reg __stream_max_pool_serial_27_stream_ivalid_5;
  reg [32-1:0] _counter_data_884;
  reg [32-1:0] _counter_count_884;
  wire _counter_reset_cond_884;
  assign _counter_reset_cond_884 = stream_max_pool_serial_27__reduce_reset_data;
  wire [32-1:0] _counter_current_count_884;
  assign _counter_current_count_884 = (_counter_reset_cond_884)? 1'sd0 : _counter_count_884;
  wire [32-1:0] _reinterpretcast_src_892;
  assign _reinterpretcast_src_892 = stream_max_pool_serial_27_source_1_data;
  wire signed [32-1:0] _reinterpretcast_data_892;
  assign _reinterpretcast_data_892 = _reinterpretcast_src_892;
  reg [4-1:0] __delay_data_1123__variable_882;
  reg signed [32-1:0] __delay_data_1124_reinterpretcast_892;
  reg [1-1:0] __delay_data_1126__variable_883;
  reg [3-1:0] __delay_data_1129__variable_880;
  reg [1-1:0] _pointer_data_887;
  reg signed [32-1:0] __delay_data_1125__delay_1124_reinterpretcast_892;
  reg [1-1:0] __delay_data_1127__delay_1126__variable_883;
  reg [3-1:0] __delay_data_1130__delay_1129__variable_880;
  reg signed [33-1:0] _cond_data_894;
  reg [1-1:0] __delay_data_1128__delay_1127__delay_1126__variable_883;
  reg [3-1:0] __delay_data_1131__delay_1130__delay_1129__variable_880;
  reg [1-1:0] __variable_wdata_271;
  assign _reduce_max_13__reduce_reset_data = __variable_wdata_271;
  reg signed [32-1:0] __variable_wdata_269;
  assign _reduce_max_13_x_data = __variable_wdata_269;
  reg [32-1:0] __variable_wdata_270;
  assign _reduce_max_13_size_data = __variable_wdata_270;
  assign __reduce_max_13_is_root = ((_stream_max_pool_serial_27_busy)? 0 : 1) && 1;
  assign __reduce_max_13_stream_oready = ((_stream_max_pool_serial_27_busy)? _stream_max_pool_serial_27_stream_oready : 1) && __reduce_max_13_stream_internal_oready;
  assign _stream_max_pool_serial_27_stream_internal_oready = ((_stream_max_pool_serial_27_busy)? __reduce_max_13_stream_internal_oready : 1) && 1;
  wire signed [32-1:0] __substreamoutput_data_896;
  assign __substreamoutput_data_896 = _reduce_max_13_data_data;
  wire [1-1:0] __substreamoutput_data_897;
  assign __substreamoutput_data_897 = _reduce_max_13_valid_data;
  wire signed [32-1:0] _reinterpretcast_src_898;
  assign _reinterpretcast_src_898 = __substreamoutput_data_896;
  wire signed [32-1:0] _reinterpretcast_data_898;
  assign _reinterpretcast_data_898 = _reinterpretcast_src_898;
  wire [1-1:0] stream_max_pool_serial_27_sink_6_data;
  assign stream_max_pool_serial_27_sink_6_data = __substreamoutput_data_897;
  wire signed [32-1:0] stream_max_pool_serial_27_sink_5_data;
  assign stream_max_pool_serial_27_sink_5_data = _reinterpretcast_data_898;
  wire _set_flag_966;
  assign _set_flag_966 = max_pool_serial_27_comp_fsm == 4;
  reg [3-1:0] __variable_wdata_880;
  assign stream_max_pool_serial_27_parameter_0_data = __variable_wdata_880;
  wire _set_flag_967;
  assign _set_flag_967 = max_pool_serial_27_comp_fsm == 4;
  reg [4-1:0] __variable_wdata_882;
  assign stream_max_pool_serial_27_parameter_2_data = __variable_wdata_882;
  reg [32-1:0] _source_stream_max_pool_serial_27_source_1_pat_cur_offset_0;
  reg [32-1:0] _source_stream_max_pool_serial_27_source_1_pat_cur_offset_1;
  reg [32-1:0] _source_stream_max_pool_serial_27_source_1_pat_cur_offset_2;
  reg [32-1:0] _source_stream_max_pool_serial_27_source_1_pat_cur_offset_3;
  reg [33-1:0] _source_stream_max_pool_serial_27_source_1_pat_size_0;
  reg [33-1:0] _source_stream_max_pool_serial_27_source_1_pat_size_1;
  reg [33-1:0] _source_stream_max_pool_serial_27_source_1_pat_size_2;
  reg [33-1:0] _source_stream_max_pool_serial_27_source_1_pat_size_3;
  reg [32-1:0] _source_stream_max_pool_serial_27_source_1_pat_stride_0;
  reg [32-1:0] _source_stream_max_pool_serial_27_source_1_pat_stride_1;
  reg [32-1:0] _source_stream_max_pool_serial_27_source_1_pat_stride_2;
  reg [32-1:0] _source_stream_max_pool_serial_27_source_1_pat_stride_3;
  reg [33-1:0] _source_stream_max_pool_serial_27_source_1_pat_count_0;
  reg [33-1:0] _source_stream_max_pool_serial_27_source_1_pat_count_1;
  reg [33-1:0] _source_stream_max_pool_serial_27_source_1_pat_count_2;
  reg [33-1:0] _source_stream_max_pool_serial_27_source_1_pat_count_3;
  reg [33-1:0] _source_stream_max_pool_serial_27_source_1_pat_size_buf_0;
  reg [33-1:0] _source_stream_max_pool_serial_27_source_1_pat_size_buf_1;
  reg [33-1:0] _source_stream_max_pool_serial_27_source_1_pat_size_buf_2;
  reg [33-1:0] _source_stream_max_pool_serial_27_source_1_pat_size_buf_3;
  reg [32-1:0] _source_stream_max_pool_serial_27_source_1_pat_stride_buf_0;
  reg [32-1:0] _source_stream_max_pool_serial_27_source_1_pat_stride_buf_1;
  reg [32-1:0] _source_stream_max_pool_serial_27_source_1_pat_stride_buf_2;
  reg [32-1:0] _source_stream_max_pool_serial_27_source_1_pat_stride_buf_3;
  wire _set_flag_968;
  assign _set_flag_968 = max_pool_serial_27_comp_fsm == 4;
  assign ram_w32_l32768_id0_0_addr = (_stream_max_pool_serial_27_stream_oready && _stream_max_pool_serial_27_source_1_source_ram_renable && (_stream_max_pool_serial_27_source_1_source_sel == 1))? _stream_max_pool_serial_27_source_1_source_ram_raddr : 'hx;
  assign ram_w32_l32768_id0_0_enable = (_stream_max_pool_serial_27_stream_oready && _stream_max_pool_serial_27_source_1_source_ram_renable && (_stream_max_pool_serial_27_source_1_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_969 = 1;
  wire [_tmp_969-1:0] _tmp_970;
  assign _tmp_970 = _stream_max_pool_serial_27_stream_oready && _stream_max_pool_serial_27_source_1_source_ram_renable && (_stream_max_pool_serial_27_source_1_source_sel == 1);
  reg [_tmp_969-1:0] __tmp_970_1;
  assign _stream_max_pool_serial_27_source_1_source_ram_rdata = (_stream_max_pool_serial_27_source_1_source_sel == 1)? ram_w32_l32768_id0_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_881;
  assign stream_max_pool_serial_27_source_1_data = __variable_wdata_881;
  reg [32-1:0] _stream_max_pool_serial_27_source_1_source_pat_fsm_0;
  localparam _stream_max_pool_serial_27_source_1_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_max_pool_serial_27_source_1_source_pat_all_offset;
  assign _stream_max_pool_serial_27_source_1_source_pat_all_offset = _stream_max_pool_serial_27_source_1_source_offset_buf + _source_stream_max_pool_serial_27_source_1_pat_cur_offset_0 + _source_stream_max_pool_serial_27_source_1_pat_cur_offset_1 + _source_stream_max_pool_serial_27_source_1_pat_cur_offset_2 + _source_stream_max_pool_serial_27_source_1_pat_cur_offset_3;
  wire _set_flag_971;
  assign _set_flag_971 = max_pool_serial_27_comp_fsm == 4;
  reg _tmp_972;
  reg _tmp_973;
  reg _tmp_974;
  reg _tmp_975;
  reg _tmp_976;
  reg _tmp_977;
  reg _tmp_978;
  localparam _tmp_979 = 33;
  wire [_tmp_979-1:0] _tmp_980;
  assign _tmp_980 = max_pool_serial_27_stream_out_local + max_pool_serial_27_out_page_comp_offset_buf;
  reg [_tmp_979-1:0] _tmp_981;
  reg [_tmp_979-1:0] _tmp_982;
  reg [_tmp_979-1:0] _tmp_983;
  reg [_tmp_979-1:0] _tmp_984;
  reg [_tmp_979-1:0] _tmp_985;
  reg [_tmp_979-1:0] _tmp_986;
  reg [_tmp_979-1:0] _tmp_987;
  reg [9-1:0] _tmp_988;
  reg [9-1:0] _tmp_989;
  reg [9-1:0] _tmp_990;
  reg [9-1:0] _tmp_991;
  reg [9-1:0] _tmp_992;
  reg [9-1:0] _tmp_993;
  reg [9-1:0] _tmp_994;
  assign ram_w32_l8192_id0_0_wdata = (_stream_max_pool_serial_27_stream_oready && _stream_max_pool_serial_27_sink_5_sink_wenable && (_stream_max_pool_serial_27_sink_5_sink_sel == 2))? _stream_max_pool_serial_27_sink_5_sink_wdata : 'hx;
  assign ram_w32_l8192_id0_0_wenable = (_stream_max_pool_serial_27_stream_oready && _stream_max_pool_serial_27_sink_5_sink_wenable && (_stream_max_pool_serial_27_sink_5_sink_sel == 2))? 1'd1 : 0;
  reg [32-1:0] _stream_max_pool_serial_27_sink_5_sink_fsm_1;
  localparam _stream_max_pool_serial_27_sink_5_sink_fsm_1_init = 0;
  wire _set_flag_995;
  assign _set_flag_995 = max_pool_serial_27_comp_fsm == 5;
  assign _stream_max_pool_serial_27_run_flag = (_set_flag_995)? 1 : 0;
  reg _tmp_996;
  reg _tmp_997;
  reg _tmp_998;
  reg _tmp_999;
  reg _tmp_1000;
  reg _tmp_1001;
  reg _tmp_1002;
  reg _tmp_1003;
  reg _tmp_1004;
  reg _tmp_1005;
  assign __reduce_max_13_source_stop = __reduce_max_13_stream_oready && 1'd0;
  reg _tmp_1006;
  reg _tmp_1007;
  reg _tmp_1008;
  assign __reduce_max_13_sink_start = _tmp_1008;
  reg _tmp_1009;
  reg _tmp_1010;
  reg _tmp_1011;
  assign __reduce_max_13_sink_stop = _tmp_1011;
  reg _tmp_1012;
  reg _tmp_1013;
  reg _tmp_1014;
  assign __reduce_max_13_sink_busy = _tmp_1014;
  reg _tmp_1015;
  assign __reduce_max_13_busy = __reduce_max_13_source_busy || __reduce_max_13_sink_busy || __reduce_max_13_busy_reg;
  reg _tmp_1016;
  reg _tmp_1017;
  reg _tmp_1018;
  reg _tmp_1019;
  reg _tmp_1020;
  reg _tmp_1021;
  reg [1-1:0] __variable_wdata_883;
  assign stream_max_pool_serial_27__reduce_reset_data = __variable_wdata_883;
  reg _tmp_1022;
  reg _tmp_1023;
  reg _tmp_1024;
  reg _tmp_1025;
  assign _stream_max_pool_serial_27_source_stop = _stream_max_pool_serial_27_stream_oready && (_stream_max_pool_serial_27_source_1_idle && (_stream_max_pool_serial_27_fsm == 3));
  localparam _tmp_1026 = 1;
  wire [_tmp_1026-1:0] _tmp_1027;
  assign _tmp_1027 = _stream_max_pool_serial_27_source_1_idle && (_stream_max_pool_serial_27_fsm == 3);
  reg [_tmp_1026-1:0] _tmp_1028;
  localparam _tmp_1029 = 1;
  wire [_tmp_1029-1:0] _tmp_1030;
  assign _tmp_1030 = _stream_max_pool_serial_27_source_1_idle && (_stream_max_pool_serial_27_fsm == 3);
  reg [_tmp_1029-1:0] _tmp_1031;
  reg _tmp_1032;
  reg _tmp_1033;
  reg _tmp_1034;
  reg _tmp_1035;
  reg _tmp_1036;
  reg _tmp_1037;
  reg _tmp_1038;
  assign _stream_max_pool_serial_27_sink_start = _tmp_1038;
  reg _tmp_1039;
  reg _tmp_1040;
  reg _tmp_1041;
  reg _tmp_1042;
  reg _tmp_1043;
  reg _tmp_1044;
  reg _tmp_1045;
  assign _stream_max_pool_serial_27_sink_stop = _tmp_1045;
  reg _tmp_1046;
  reg _tmp_1047;
  reg _tmp_1048;
  reg _tmp_1049;
  reg _tmp_1050;
  reg _tmp_1051;
  reg _tmp_1052;
  assign _stream_max_pool_serial_27_sink_busy = _tmp_1052;
  reg _tmp_1053;
  assign _stream_max_pool_serial_27_busy = _stream_max_pool_serial_27_source_busy || _stream_max_pool_serial_27_sink_busy || _stream_max_pool_serial_27_busy_reg;
  wire [32-1:0] mask_addr_shifted_1054;
  assign mask_addr_shifted_1054 = max_pool_serial_27_objaddr + max_pool_serial_27_out_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1055;
  assign mask_addr_masked_1055 = mask_addr_shifted_1054 << 2;
  reg [32-1:0] read_burst_fsm_26;
  localparam read_burst_fsm_26_init = 0;
  reg [13-1:0] read_burst_addr_1056;
  reg [13-1:0] read_burst_stride_1057;
  reg [33-1:0] read_burst_length_1058;
  reg read_burst_rvalid_1059;
  reg read_burst_rlast_1060;
  localparam _tmp_1061 = 1;
  wire [_tmp_1061-1:0] _tmp_1062;
  assign _tmp_1062 = (read_burst_fsm_26 == 1) && (!read_burst_rvalid_1059 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1061-1:0] __tmp_1062_1;
  wire [32-1:0] read_burst_rdata_1063;
  assign read_burst_rdata_1063 = ram_w32_l8192_id0_1_rdata;
  reg _maxi_wdata_cond_1_1;
  reg [32-1:0] max_pool_47_objaddr;
  reg [32-1:0] max_pool_47_arg_objaddr_0;
  reg [32-1:0] control_max_pool_47;
  localparam control_max_pool_47_init = 0;
  reg _control_max_pool_47_called;
  wire signed [32-1:0] max_pool_47_act_base_offset;
  reg signed [32-1:0] max_pool_47_act_base_offset_row;
  reg signed [32-1:0] max_pool_47_act_base_offset_bat;
  assign max_pool_47_act_base_offset = max_pool_47_act_base_offset_row + max_pool_47_act_base_offset_bat;
  wire signed [32-1:0] max_pool_47_out_base_offset;
  reg signed [32-1:0] max_pool_47_out_base_offset_row;
  reg signed [32-1:0] max_pool_47_out_base_offset_bat;
  assign max_pool_47_out_base_offset = max_pool_47_out_base_offset_row + max_pool_47_out_base_offset_bat;
  reg max_pool_47_dma_flag_0;
  reg max_pool_47_dma_flag_1;
  reg [32-1:0] max_pool_47_col_count;
  reg [32-1:0] max_pool_47_row_count;
  reg [32-1:0] max_pool_47_bat_count;
  reg [1-1:0] max_pool_47_col_select;
  reg [1-1:0] max_pool_47_row_select;
  reg [32-1:0] max_pool_47_prev_row_count;
  reg [32-1:0] max_pool_47_prev_bat_count;
  reg [1-1:0] max_pool_47_prev_row_select;
  reg [32-1:0] max_pool_47_stream_act_local_0;
  reg [32-1:0] max_pool_47_stream_act_local_1;
  reg [32-1:0] max_pool_47_stream_act_local_2;
  reg [32-1:0] max_pool_47_stream_act_local_3;
  reg [32-1:0] max_pool_47_stream_out_local;
  reg max_pool_47_act_page_0;
  reg max_pool_47_act_page_1;
  reg [32-1:0] max_pool_47_act_page_comp_offset_0;
  reg [32-1:0] max_pool_47_act_page_comp_offset_1;
  reg [32-1:0] max_pool_47_act_page_dma_offset_0;
  reg [32-1:0] max_pool_47_act_page_dma_offset_1;
  reg max_pool_47_out_page;
  reg [32-1:0] max_pool_47_out_page_comp_offset;
  reg [32-1:0] max_pool_47_out_page_dma_offset;
  reg max_pool_47_skip_read_act;
  reg max_pool_47_skip_comp;
  reg max_pool_47_skip_write_out;
  reg [32-1:0] max_pool_47_comp_count;
  reg [32-1:0] max_pool_47_out_count;
  wire max_pool_47_dma_pad_mask_0;
  assign max_pool_47_dma_pad_mask_0 = (max_pool_47_row_count + 0 < cparam_max_pool_47_pad_row_top) || (max_pool_47_row_count + 0 >= cparam_max_pool_47_act_num_row + cparam_max_pool_47_pad_row_top);
  wire max_pool_47_dma_pad_mask_1;
  assign max_pool_47_dma_pad_mask_1 = (max_pool_47_row_count + 1 < cparam_max_pool_47_pad_row_top) || (max_pool_47_row_count + 1 >= cparam_max_pool_47_act_num_row + cparam_max_pool_47_pad_row_top);
  wire [32-1:0] max_pool_47_mux_act_gaddr_0;
  assign max_pool_47_mux_act_gaddr_0 = (max_pool_47_row_select == 0)? max_pool_47_arg_objaddr_0 + (max_pool_47_act_base_offset + cparam_max_pool_47_act_offset_values_0) : 
                                       (max_pool_47_row_select == 1)? max_pool_47_arg_objaddr_0 + (max_pool_47_act_base_offset + cparam_max_pool_47_act_offset_values_1) : 1'd0;
  wire [32-1:0] max_pool_47_mux_act_gaddr_1;
  assign max_pool_47_mux_act_gaddr_1 = (max_pool_47_row_select == 0)? max_pool_47_arg_objaddr_0 + (max_pool_47_act_base_offset + cparam_max_pool_47_act_offset_values_1) : 
                                       (max_pool_47_row_select == 1)? max_pool_47_arg_objaddr_0 + (max_pool_47_act_base_offset + cparam_max_pool_47_act_offset_values_0) : 1'd0;
  wire max_pool_47_mux_dma_pad_mask_0;
  assign max_pool_47_mux_dma_pad_mask_0 = (max_pool_47_row_select == 0)? max_pool_47_dma_pad_mask_0 : 
                                          (max_pool_47_row_select == 1)? max_pool_47_dma_pad_mask_1 : 1'd0;
  wire max_pool_47_mux_dma_pad_mask_1;
  assign max_pool_47_mux_dma_pad_mask_1 = (max_pool_47_row_select == 0)? max_pool_47_dma_pad_mask_1 : 
                                          (max_pool_47_row_select == 1)? max_pool_47_dma_pad_mask_0 : 1'd0;
  wire max_pool_47_mux_dma_flag_0;
  assign max_pool_47_mux_dma_flag_0 = (max_pool_47_prev_row_select == 0)? max_pool_47_dma_flag_0 : 
                                      (max_pool_47_prev_row_select == 1)? max_pool_47_dma_flag_1 : 1'd0;
  wire max_pool_47_mux_dma_flag_1;
  assign max_pool_47_mux_dma_flag_1 = (max_pool_47_prev_row_select == 0)? max_pool_47_dma_flag_1 : 
                                      (max_pool_47_prev_row_select == 1)? max_pool_47_dma_flag_0 : 1'd0;
  wire [32-1:0] mask_addr_shifted_1064;
  assign mask_addr_shifted_1064 = max_pool_47_mux_act_gaddr_0 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1065;
  assign mask_addr_masked_1065 = mask_addr_shifted_1064 << 2;
  wire write_burst_block_ram_wvalid_1066;
  wire write_burst_block_ram_wquit_1067;
  reg [32-1:0] write_burst_fsm_27;
  localparam write_burst_fsm_27_init = 0;
  reg [13-1:0] write_burst_addr_1068;
  reg [13-1:0] write_burst_stride_1069;
  reg [33-1:0] write_burst_length_1070;
  reg write_burst_done_1071;
  assign ram_w32_l8192_id0_1_addr = ((write_burst_fsm_27 == 1) && write_burst_block_ram_wvalid_1066)? write_burst_addr_1068 : 
                                    ((read_burst_fsm_26 == 1) && (!read_burst_rvalid_1059 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_addr_1056 : 
                                    ((write_burst_fsm_22 == 1) && write_burst_block_ram_wvalid_208)? write_burst_addr_210 : 'hx;
  assign ram_w32_l8192_id0_1_wdata = ((write_burst_fsm_27 == 1) && write_burst_block_ram_wvalid_1066)? _maxi_rdata_sb_0 : 
                                     ((write_burst_fsm_22 == 1) && write_burst_block_ram_wvalid_208)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l8192_id0_1_wenable = ((write_burst_fsm_27 == 1) && write_burst_block_ram_wvalid_1066)? 1'd1 : 
                                       ((write_burst_fsm_22 == 1) && write_burst_block_ram_wvalid_208)? 1'd1 : 0;
  assign ram_w32_l8192_id0_1_enable = ((write_burst_fsm_27 == 1) && write_burst_block_ram_wvalid_1066)? 1'd1 : 
                                      ((read_burst_fsm_26 == 1) && (!read_burst_rvalid_1059 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 
                                      ((write_burst_fsm_22 == 1) && write_burst_block_ram_wvalid_208)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_1072;
  wire write_burst_block_ram_wquit_1073;
  reg [32-1:0] write_burst_fsm_28;
  localparam write_burst_fsm_28_init = 0;
  reg [13-1:0] write_burst_addr_1074;
  reg [13-1:0] write_burst_stride_1075;
  reg [33-1:0] write_burst_length_1076;
  reg write_burst_done_1077;
  assign ram_w32_l8192_id1_1_addr = ((write_burst_fsm_28 == 1) && write_burst_block_ram_wvalid_1072)? write_burst_addr_1074 : 'hx;
  assign ram_w32_l8192_id1_1_wdata = ((write_burst_fsm_28 == 1) && write_burst_block_ram_wvalid_1072)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l8192_id1_1_wenable = ((write_burst_fsm_28 == 1) && write_burst_block_ram_wvalid_1072)? 1'd1 : 0;
  assign ram_w32_l8192_id1_1_enable = ((write_burst_fsm_28 == 1) && write_burst_block_ram_wvalid_1072)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_29;
  localparam write_burst_block_fsm_29_init = 0;
  reg [33-1:0] write_burst_block_length_1078;
  reg [32-1:0] write_burst_block_blocksize_1079;
  reg write_burst_block_done_1080;
  reg [32-1:0] write_burst_block_count_1081;
  assign write_burst_block_ram_wvalid_1066 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_29 == 1);
  assign write_burst_block_ram_wquit_1067 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_1078 <= 1);
  assign write_burst_block_ram_wvalid_1072 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_29 == 2);
  assign write_burst_block_ram_wquit_1073 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_1078 <= 1);
  wire [32-1:0] mask_addr_shifted_1082;
  assign mask_addr_shifted_1082 = max_pool_47_mux_act_gaddr_1 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1083;
  assign mask_addr_masked_1083 = mask_addr_shifted_1082 << 2;
  assign _maxi_read_req_fifo_deq = ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 9)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 8)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 7)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 6)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1)) && !_maxi_read_req_fifo_empty)? 1 : 0;
  wire write_burst_block_ram_wvalid_1084;
  wire write_burst_block_ram_wquit_1085;
  reg [32-1:0] write_burst_fsm_30;
  localparam write_burst_fsm_30_init = 0;
  reg [13-1:0] write_burst_addr_1086;
  reg [13-1:0] write_burst_stride_1087;
  reg [33-1:0] write_burst_length_1088;
  reg write_burst_done_1089;
  assign ram_w32_l8192_id2_1_addr = ((write_burst_fsm_30 == 1) && write_burst_block_ram_wvalid_1084)? write_burst_addr_1086 : 'hx;
  assign ram_w32_l8192_id2_1_wdata = ((write_burst_fsm_30 == 1) && write_burst_block_ram_wvalid_1084)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l8192_id2_1_wenable = ((write_burst_fsm_30 == 1) && write_burst_block_ram_wvalid_1084)? 1'd1 : 0;
  assign ram_w32_l8192_id2_1_enable = ((write_burst_fsm_30 == 1) && write_burst_block_ram_wvalid_1084)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_1090;
  wire write_burst_block_ram_wquit_1091;
  reg [32-1:0] write_burst_fsm_31;
  localparam write_burst_fsm_31_init = 0;
  reg [13-1:0] write_burst_addr_1092;
  reg [13-1:0] write_burst_stride_1093;
  reg [33-1:0] write_burst_length_1094;
  reg write_burst_done_1095;
  assign ram_w32_l8192_id3_1_addr = ((write_burst_fsm_31 == 1) && write_burst_block_ram_wvalid_1090)? write_burst_addr_1092 : 'hx;
  assign ram_w32_l8192_id3_1_wdata = ((write_burst_fsm_31 == 1) && write_burst_block_ram_wvalid_1090)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l8192_id3_1_wenable = ((write_burst_fsm_31 == 1) && write_burst_block_ram_wvalid_1090)? 1'd1 : 0;
  assign ram_w32_l8192_id3_1_enable = ((write_burst_fsm_31 == 1) && write_burst_block_ram_wvalid_1090)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_32;
  localparam write_burst_block_fsm_32_init = 0;
  reg [33-1:0] write_burst_block_length_1096;
  reg [32-1:0] write_burst_block_blocksize_1097;
  reg write_burst_block_done_1098;
  reg [32-1:0] write_burst_block_count_1099;
  assign write_burst_block_ram_wvalid_1084 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_32 == 1);
  assign write_burst_block_ram_wquit_1085 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_1096 <= 1);
  assign write_burst_block_ram_wvalid_1090 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_32 == 2);
  assign write_burst_block_ram_wquit_1091 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_1096 <= 1);
  assign _maxi_rready_sb_0 = (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2);
  reg [32-1:0] max_pool_47_comp_fsm;
  localparam max_pool_47_comp_fsm_init = 0;
  reg [32-1:0] max_pool_47_act_page_comp_offset_buf_0;
  reg [32-1:0] max_pool_47_act_page_comp_offset_buf_1;
  reg [32-1:0] max_pool_47_out_page_comp_offset_buf;
  reg [32-1:0] max_pool_47_row_count_buf;
  reg [1-1:0] max_pool_47_row_select_buf;
  wire max_pool_47_stream_pad_mask_0_0;
  assign max_pool_47_stream_pad_mask_0_0 = (max_pool_47_col_count + 0 < cparam_max_pool_47_pad_col_left) || (max_pool_47_col_count + 0 >= cparam_max_pool_47_act_num_col + cparam_max_pool_47_pad_col_left) || (max_pool_47_row_count_buf + 0 < cparam_max_pool_47_pad_row_top) || (max_pool_47_row_count_buf + 0 >= cparam_max_pool_47_act_num_row + cparam_max_pool_47_pad_row_top);
  wire max_pool_47_stream_pad_mask_0_1;
  assign max_pool_47_stream_pad_mask_0_1 = (max_pool_47_col_count + 1 < cparam_max_pool_47_pad_col_left) || (max_pool_47_col_count + 1 >= cparam_max_pool_47_act_num_col + cparam_max_pool_47_pad_col_left) || (max_pool_47_row_count_buf + 0 < cparam_max_pool_47_pad_row_top) || (max_pool_47_row_count_buf + 0 >= cparam_max_pool_47_act_num_row + cparam_max_pool_47_pad_row_top);
  wire max_pool_47_stream_pad_mask_1_0;
  assign max_pool_47_stream_pad_mask_1_0 = (max_pool_47_col_count + 0 < cparam_max_pool_47_pad_col_left) || (max_pool_47_col_count + 0 >= cparam_max_pool_47_act_num_col + cparam_max_pool_47_pad_col_left) || (max_pool_47_row_count_buf + 1 < cparam_max_pool_47_pad_row_top) || (max_pool_47_row_count_buf + 1 >= cparam_max_pool_47_act_num_row + cparam_max_pool_47_pad_row_top);
  wire max_pool_47_stream_pad_mask_1_1;
  assign max_pool_47_stream_pad_mask_1_1 = (max_pool_47_col_count + 1 < cparam_max_pool_47_pad_col_left) || (max_pool_47_col_count + 1 >= cparam_max_pool_47_act_num_col + cparam_max_pool_47_pad_col_left) || (max_pool_47_row_count_buf + 1 < cparam_max_pool_47_pad_row_top) || (max_pool_47_row_count_buf + 1 >= cparam_max_pool_47_act_num_row + cparam_max_pool_47_pad_row_top);
  reg [4-1:0] max_pool_47_stream_pad_masks;
  wire [4-1:0] stream_max_pool_47_parameter_0_data;
  wire [32-1:0] stream_max_pool_47_source_1_data;
  wire [32-1:0] stream_max_pool_47_source_2_data;
  wire [32-1:0] stream_max_pool_47_source_3_data;
  wire [32-1:0] stream_max_pool_47_source_4_data;
  reg __stream_max_pool_47_stream_ivalid_1;
  reg __stream_max_pool_47_stream_ivalid_2;
  reg __stream_max_pool_47_stream_ivalid_3;
  reg __stream_max_pool_47_stream_ivalid_4;
  reg __stream_max_pool_47_stream_ivalid_5;
  reg __stream_max_pool_47_stream_ivalid_6;
  wire [32-1:0] _reinterpretcast_src_920;
  assign _reinterpretcast_src_920 = stream_max_pool_47_source_1_data;
  wire signed [32-1:0] _reinterpretcast_data_920;
  assign _reinterpretcast_data_920 = _reinterpretcast_src_920;
  wire [32-1:0] _reinterpretcast_src_921;
  assign _reinterpretcast_src_921 = stream_max_pool_47_source_2_data;
  wire signed [32-1:0] _reinterpretcast_data_921;
  assign _reinterpretcast_data_921 = _reinterpretcast_src_921;
  wire [32-1:0] _reinterpretcast_src_922;
  assign _reinterpretcast_src_922 = stream_max_pool_47_source_3_data;
  wire signed [32-1:0] _reinterpretcast_data_922;
  assign _reinterpretcast_data_922 = _reinterpretcast_src_922;
  wire [32-1:0] _reinterpretcast_src_923;
  assign _reinterpretcast_src_923 = stream_max_pool_47_source_4_data;
  wire signed [32-1:0] _reinterpretcast_data_923;
  assign _reinterpretcast_data_923 = _reinterpretcast_src_923;
  wire [1-1:0] _pointer_data_925;
  assign _pointer_data_925 = stream_max_pool_47_parameter_0_data[1'sd0];
  reg signed [33-1:0] _cond_data_927;
  wire [1-1:0] _pointer_data_928;
  assign _pointer_data_928 = stream_max_pool_47_parameter_0_data[2'sd1];
  reg signed [33-1:0] _cond_data_930;
  wire [1-1:0] _pointer_data_931;
  assign _pointer_data_931 = stream_max_pool_47_parameter_0_data[3'sd2];
  reg signed [33-1:0] _cond_data_933;
  wire [1-1:0] _pointer_data_934;
  assign _pointer_data_934 = stream_max_pool_47_parameter_0_data[3'sd3];
  reg signed [33-1:0] _cond_data_936;
  reg signed [32-1:0] __variable_wdata_0;
  assign _max_0_var0_data = __variable_wdata_0;
  reg signed [32-1:0] __variable_wdata_1;
  assign _max_0_var1_data = __variable_wdata_1;
  reg signed [32-1:0] __variable_wdata_2;
  assign _max_0_var2_data = __variable_wdata_2;
  reg signed [32-1:0] __variable_wdata_3;
  assign _max_0_var3_data = __variable_wdata_3;
  assign __max_0_is_root = ((_stream_max_pool_47_busy)? 0 : 1) && 1;
  assign __max_0_stream_oready = ((_stream_max_pool_47_busy)? _stream_max_pool_47_stream_oready : 1) && __max_0_stream_internal_oready;
  assign _stream_max_pool_47_stream_internal_oready = ((_stream_max_pool_47_busy)? __max_0_stream_internal_oready : 1) && 1;
  wire signed [32-1:0] __substreamoutput_data_944;
  assign __substreamoutput_data_944 = _max_0_val_data;
  wire signed [32-1:0] _reinterpretcast_src_945;
  assign _reinterpretcast_src_945 = __substreamoutput_data_944;
  wire signed [32-1:0] _reinterpretcast_data_945;
  assign _reinterpretcast_data_945 = _reinterpretcast_src_945;
  wire signed [32-1:0] stream_max_pool_47_sink_6_data;
  assign stream_max_pool_47_sink_6_data = _reinterpretcast_data_945;
  wire _set_flag_1100;
  assign _set_flag_1100 = max_pool_47_comp_fsm == 4;
  reg [4-1:0] __variable_wdata_899;
  assign stream_max_pool_47_parameter_0_data = __variable_wdata_899;
  wire _set_flag_1101;
  assign _set_flag_1101 = max_pool_47_comp_fsm == 4;
  assign ram_w32_l8192_id0_0_addr = (_stream_max_pool_47_stream_oready && _stream_max_pool_47_source_1_source_ram_renable && (_stream_max_pool_47_source_1_source_sel == 1))? _stream_max_pool_47_source_1_source_ram_raddr : 
                                    (_stream_max_pool_serial_27_stream_oready && _stream_max_pool_serial_27_sink_5_sink_wenable && (_stream_max_pool_serial_27_sink_5_sink_sel == 2))? _stream_max_pool_serial_27_sink_5_sink_waddr : 
                                    (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_28_source_ram_renable && (_stream_conv2d_25_source_28_source_sel == 11))? _stream_conv2d_25_source_28_source_ram_raddr : 'hx;
  assign ram_w32_l8192_id0_0_enable = (_stream_max_pool_47_stream_oready && _stream_max_pool_47_source_1_source_ram_renable && (_stream_max_pool_47_source_1_source_sel == 1))? 1'd1 : 
                                      (_stream_max_pool_serial_27_stream_oready && _stream_max_pool_serial_27_sink_5_sink_wenable && (_stream_max_pool_serial_27_sink_5_sink_sel == 2))? 1'd1 : 
                                      (_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_28_source_ram_renable && (_stream_conv2d_25_source_28_source_sel == 11))? 1'd1 : 0;
  localparam _tmp_1102 = 1;
  wire [_tmp_1102-1:0] _tmp_1103;
  assign _tmp_1103 = _stream_max_pool_47_stream_oready && _stream_max_pool_47_source_1_source_ram_renable && (_stream_max_pool_47_source_1_source_sel == 1);
  reg [_tmp_1102-1:0] __tmp_1103_1;
  assign _stream_max_pool_47_source_1_source_ram_rdata = (_stream_max_pool_47_source_1_source_sel == 1)? ram_w32_l8192_id0_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_900;
  assign stream_max_pool_47_source_1_data = __variable_wdata_900;
  reg [32-1:0] _stream_max_pool_47_source_1_source_fsm_0;
  localparam _stream_max_pool_47_source_1_source_fsm_0_init = 0;
  wire _set_flag_1104;
  assign _set_flag_1104 = max_pool_47_comp_fsm == 4;
  assign ram_w32_l8192_id1_0_addr = (_stream_max_pool_47_stream_oready && _stream_max_pool_47_source_2_source_ram_renable && (_stream_max_pool_47_source_2_source_sel == 2))? _stream_max_pool_47_source_2_source_ram_raddr : 'hx;
  assign ram_w32_l8192_id1_0_enable = (_stream_max_pool_47_stream_oready && _stream_max_pool_47_source_2_source_ram_renable && (_stream_max_pool_47_source_2_source_sel == 2))? 1'd1 : 0;
  localparam _tmp_1105 = 1;
  wire [_tmp_1105-1:0] _tmp_1106;
  assign _tmp_1106 = _stream_max_pool_47_stream_oready && _stream_max_pool_47_source_2_source_ram_renable && (_stream_max_pool_47_source_2_source_sel == 2);
  reg [_tmp_1105-1:0] __tmp_1106_1;
  assign _stream_max_pool_47_source_2_source_ram_rdata = (_stream_max_pool_47_source_2_source_sel == 2)? ram_w32_l8192_id1_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_901;
  assign stream_max_pool_47_source_2_data = __variable_wdata_901;
  reg [32-1:0] _stream_max_pool_47_source_2_source_fsm_1;
  localparam _stream_max_pool_47_source_2_source_fsm_1_init = 0;
  wire _set_flag_1107;
  assign _set_flag_1107 = max_pool_47_comp_fsm == 4;
  assign ram_w32_l8192_id2_0_addr = (_stream_max_pool_47_stream_oready && _stream_max_pool_47_source_3_source_ram_renable && (_stream_max_pool_47_source_3_source_sel == 3))? _stream_max_pool_47_source_3_source_ram_raddr : 'hx;
  assign ram_w32_l8192_id2_0_enable = (_stream_max_pool_47_stream_oready && _stream_max_pool_47_source_3_source_ram_renable && (_stream_max_pool_47_source_3_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_1108 = 1;
  wire [_tmp_1108-1:0] _tmp_1109;
  assign _tmp_1109 = _stream_max_pool_47_stream_oready && _stream_max_pool_47_source_3_source_ram_renable && (_stream_max_pool_47_source_3_source_sel == 3);
  reg [_tmp_1108-1:0] __tmp_1109_1;
  assign _stream_max_pool_47_source_3_source_ram_rdata = (_stream_max_pool_47_source_3_source_sel == 3)? ram_w32_l8192_id2_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_902;
  assign stream_max_pool_47_source_3_data = __variable_wdata_902;
  reg [32-1:0] _stream_max_pool_47_source_3_source_fsm_2;
  localparam _stream_max_pool_47_source_3_source_fsm_2_init = 0;
  wire _set_flag_1110;
  assign _set_flag_1110 = max_pool_47_comp_fsm == 4;
  assign ram_w32_l8192_id3_0_addr = (_stream_max_pool_47_stream_oready && _stream_max_pool_47_source_4_source_ram_renable && (_stream_max_pool_47_source_4_source_sel == 4))? _stream_max_pool_47_source_4_source_ram_raddr : 'hx;
  assign ram_w32_l8192_id3_0_enable = (_stream_max_pool_47_stream_oready && _stream_max_pool_47_source_4_source_ram_renable && (_stream_max_pool_47_source_4_source_sel == 4))? 1'd1 : 0;
  localparam _tmp_1111 = 1;
  wire [_tmp_1111-1:0] _tmp_1112;
  assign _tmp_1112 = _stream_max_pool_47_stream_oready && _stream_max_pool_47_source_4_source_ram_renable && (_stream_max_pool_47_source_4_source_sel == 4);
  reg [_tmp_1111-1:0] __tmp_1112_1;
  assign _stream_max_pool_47_source_4_source_ram_rdata = (_stream_max_pool_47_source_4_source_sel == 4)? ram_w32_l8192_id3_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_903;
  assign stream_max_pool_47_source_4_data = __variable_wdata_903;
  reg [32-1:0] _stream_max_pool_47_source_4_source_fsm_3;
  localparam _stream_max_pool_47_source_4_source_fsm_3_init = 0;
  wire _set_flag_1113;
  assign _set_flag_1113 = max_pool_47_comp_fsm == 4;
  reg _tmp_1114;
  reg _tmp_1115;
  reg _tmp_1116;
  reg _tmp_1117;
  reg _tmp_1118;
  reg _tmp_1119;
  reg _tmp_1120;
  reg _tmp_1121;
  localparam _tmp_1122 = 33;
  wire [_tmp_1122-1:0] _tmp_1123;
  assign _tmp_1123 = max_pool_47_stream_out_local + max_pool_47_out_page_comp_offset_buf;
  reg [_tmp_1122-1:0] _tmp_1124;
  reg [_tmp_1122-1:0] _tmp_1125;
  reg [_tmp_1122-1:0] _tmp_1126;
  reg [_tmp_1122-1:0] _tmp_1127;
  reg [_tmp_1122-1:0] _tmp_1128;
  reg [_tmp_1122-1:0] _tmp_1129;
  reg [_tmp_1122-1:0] _tmp_1130;
  reg [_tmp_1122-1:0] _tmp_1131;
  reg [10-1:0] _tmp_1132;
  reg [10-1:0] _tmp_1133;
  reg [10-1:0] _tmp_1134;
  reg [10-1:0] _tmp_1135;
  reg [10-1:0] _tmp_1136;
  reg [10-1:0] _tmp_1137;
  reg [10-1:0] _tmp_1138;
  reg [10-1:0] _tmp_1139;
  assign ram_w32_l16384_id0_0_addr = (_stream_max_pool_47_stream_oready && _stream_max_pool_47_sink_6_sink_wenable && (_stream_max_pool_47_sink_6_sink_sel == 5))? _stream_max_pool_47_sink_6_sink_waddr : 'hx;
  assign ram_w32_l16384_id0_0_wdata = (_stream_max_pool_47_stream_oready && _stream_max_pool_47_sink_6_sink_wenable && (_stream_max_pool_47_sink_6_sink_sel == 5))? _stream_max_pool_47_sink_6_sink_wdata : 'hx;
  assign ram_w32_l16384_id0_0_wenable = (_stream_max_pool_47_stream_oready && _stream_max_pool_47_sink_6_sink_wenable && (_stream_max_pool_47_sink_6_sink_sel == 5))? 1'd1 : 0;
  assign ram_w32_l16384_id0_0_enable = (_stream_max_pool_47_stream_oready && _stream_max_pool_47_sink_6_sink_wenable && (_stream_max_pool_47_sink_6_sink_sel == 5))? 1'd1 : 0;
  reg [32-1:0] _stream_max_pool_47_sink_6_sink_fsm_4;
  localparam _stream_max_pool_47_sink_6_sink_fsm_4_init = 0;
  wire _set_flag_1140;
  assign _set_flag_1140 = max_pool_47_comp_fsm == 5;
  assign _stream_max_pool_47_run_flag = (_set_flag_1140)? 1 : 0;
  reg _tmp_1141;
  reg _tmp_1142;
  reg _tmp_1143;
  assign __max_0_source_stop = __max_0_stream_oready && 1'd0;
  reg _tmp_1144;
  reg _tmp_1145;
  reg _tmp_1146;
  reg _tmp_1147;
  reg _tmp_1148;
  reg _tmp_1149;
  assign __max_0_sink_start = _tmp_1149;
  reg _tmp_1150;
  reg _tmp_1151;
  reg _tmp_1152;
  reg _tmp_1153;
  reg _tmp_1154;
  reg _tmp_1155;
  assign __max_0_sink_stop = _tmp_1155;
  reg _tmp_1156;
  reg _tmp_1157;
  reg _tmp_1158;
  reg _tmp_1159;
  reg _tmp_1160;
  reg _tmp_1161;
  assign __max_0_sink_busy = _tmp_1161;
  reg _tmp_1162;
  assign __max_0_busy = __max_0_source_busy || __max_0_sink_busy || __max_0_busy_reg;
  reg _tmp_1163;
  reg _tmp_1164;
  reg _tmp_1165;
  assign _stream_max_pool_47_source_stop = _stream_max_pool_47_stream_oready && (_stream_max_pool_47_source_1_idle && _stream_max_pool_47_source_2_idle && _stream_max_pool_47_source_3_idle && _stream_max_pool_47_source_4_idle && (_stream_max_pool_47_fsm == 3));
  localparam _tmp_1166 = 1;
  wire [_tmp_1166-1:0] _tmp_1167;
  assign _tmp_1167 = _stream_max_pool_47_source_1_idle && _stream_max_pool_47_source_2_idle && _stream_max_pool_47_source_3_idle && _stream_max_pool_47_source_4_idle && (_stream_max_pool_47_fsm == 3);
  reg [_tmp_1166-1:0] _tmp_1168;
  reg _tmp_1169;
  reg _tmp_1170;
  reg _tmp_1171;
  reg _tmp_1172;
  reg _tmp_1173;
  reg _tmp_1174;
  reg _tmp_1175;
  reg _tmp_1176;
  assign _stream_max_pool_47_sink_start = _tmp_1176;
  reg _tmp_1177;
  reg _tmp_1178;
  reg _tmp_1179;
  reg _tmp_1180;
  reg _tmp_1181;
  reg _tmp_1182;
  reg _tmp_1183;
  reg _tmp_1184;
  assign _stream_max_pool_47_sink_stop = _tmp_1184;
  reg _tmp_1185;
  reg _tmp_1186;
  reg _tmp_1187;
  reg _tmp_1188;
  reg _tmp_1189;
  reg _tmp_1190;
  reg _tmp_1191;
  reg _tmp_1192;
  assign _stream_max_pool_47_sink_busy = _tmp_1192;
  reg _tmp_1193;
  assign _stream_max_pool_47_busy = _stream_max_pool_47_source_busy || _stream_max_pool_47_sink_busy || _stream_max_pool_47_busy_reg;
  wire [32-1:0] mask_addr_shifted_1194;
  assign mask_addr_shifted_1194 = max_pool_47_objaddr + max_pool_47_out_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1195;
  assign mask_addr_masked_1195 = mask_addr_shifted_1194 << 2;
  reg [32-1:0] read_burst_fsm_33;
  localparam read_burst_fsm_33_init = 0;
  reg [14-1:0] read_burst_addr_1196;
  reg [14-1:0] read_burst_stride_1197;
  reg [33-1:0] read_burst_length_1198;
  reg read_burst_rvalid_1199;
  reg read_burst_rlast_1200;
  assign ram_w32_l16384_id0_1_addr = ((read_burst_fsm_33 == 1) && (!read_burst_rvalid_1199 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_addr_1196 : 'hx;
  assign ram_w32_l16384_id0_1_enable = ((read_burst_fsm_33 == 1) && (!read_burst_rvalid_1199 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 0;
  localparam _tmp_1201 = 1;
  wire [_tmp_1201-1:0] _tmp_1202;
  assign _tmp_1202 = (read_burst_fsm_33 == 1) && (!read_burst_rvalid_1199 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1201-1:0] __tmp_1202_1;
  wire [32-1:0] read_burst_rdata_1203;
  assign read_burst_rdata_1203 = ram_w32_l16384_id0_1_rdata;
  assign _maxi_write_req_fifo_deq = ((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 3)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1)) && !_maxi_write_req_fifo_empty)? 1 : 0;
  reg _maxi_wdata_cond_2_1;
  wire max_pool_47_mux_next_dma_flag_0;
  assign max_pool_47_mux_next_dma_flag_0 = (max_pool_47_row_select == 0)? (max_pool_47_row_count >= cparam_max_pool_47_max_row_count)? 1 : cparam_max_pool_47_dma_flag_conds_0 : 
                                           (max_pool_47_row_select == 1)? (max_pool_47_row_count >= cparam_max_pool_47_max_row_count)? 1 : cparam_max_pool_47_dma_flag_conds_1 : 1'd0;
  wire max_pool_47_mux_next_dma_flag_1;
  assign max_pool_47_mux_next_dma_flag_1 = (max_pool_47_row_select == 0)? (max_pool_47_row_count >= cparam_max_pool_47_max_row_count)? 1 : cparam_max_pool_47_dma_flag_conds_1 : 
                                           (max_pool_47_row_select == 1)? (max_pool_47_row_count >= cparam_max_pool_47_max_row_count)? 1 : cparam_max_pool_47_dma_flag_conds_0 : 1'd0;

  always @(posedge CLK) begin
    _RESETN_inv_1 <= RESETN_inv;
    _RESETN_inv_2 <= _RESETN_inv_1;
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      maxi_awaddr <= 0;
      maxi_awlen <= 0;
      maxi_awvalid <= 0;
      _maxi_waddr_cond_0_1 <= 0;
    end else begin
      if(_maxi_waddr_cond_0_1) begin
        maxi_awvalid <= 0;
      end 
      if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (_maxi_outstanding_wcount < 6) && ((_maxi_outstanding_wcount < 6) && (maxi_awready || !maxi_awvalid))) begin
        maxi_awaddr <= _maxi_write_global_addr;
        maxi_awlen <= _maxi_write_cur_global_size - 1;
        maxi_awvalid <= 1;
      end 
      if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (_maxi_outstanding_wcount < 6) && ((_maxi_outstanding_wcount < 6) && (maxi_awready || !maxi_awvalid)) && (_maxi_write_cur_global_size == 0)) begin
        maxi_awvalid <= 0;
      end 
      _maxi_waddr_cond_0_1 <= 1;
      if(maxi_awvalid && !maxi_awready) begin
        maxi_awvalid <= maxi_awvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_wdata_sb_0 <= 0;
      _maxi_wvalid_sb_0 <= 0;
      _maxi_wlast_sb_0 <= 0;
      _maxi_wstrb_sb_0 <= 0;
      _maxi_wdata_cond_0_1 <= 0;
      _maxi_wdata_cond_1_1 <= 0;
      _maxi_wdata_cond_2_1 <= 0;
    end else begin
      if(_maxi_wdata_cond_0_1) begin
        _maxi_wvalid_sb_0 <= 0;
        _maxi_wlast_sb_0 <= 0;
      end 
      if(_maxi_wdata_cond_1_1) begin
        _maxi_wvalid_sb_0 <= 0;
        _maxi_wlast_sb_0 <= 0;
      end 
      if(_maxi_wdata_cond_2_1) begin
        _maxi_wvalid_sb_0 <= 0;
        _maxi_wlast_sb_0 <= 0;
      end 
      if((_maxi_write_op_sel_buf == 1) && read_burst_rvalid_953 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0)) begin
        _maxi_wdata_sb_0 <= read_burst_rdata_957;
        _maxi_wvalid_sb_0 <= 1;
        _maxi_wlast_sb_0 <= read_burst_rlast_954 || (_maxi_write_size_buf == 1);
        _maxi_wstrb_sb_0 <= { 4{ 1'd1 } };
      end 
      _maxi_wdata_cond_0_1 <= 1;
      if(_maxi_wvalid_sb_0 && !_maxi_wready_sb_0) begin
        _maxi_wvalid_sb_0 <= _maxi_wvalid_sb_0;
        _maxi_wlast_sb_0 <= _maxi_wlast_sb_0;
      end 
      if((_maxi_write_op_sel_buf == 2) && read_burst_rvalid_1059 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0)) begin
        _maxi_wdata_sb_0 <= read_burst_rdata_1063;
        _maxi_wvalid_sb_0 <= 1;
        _maxi_wlast_sb_0 <= read_burst_rlast_1060 || (_maxi_write_size_buf == 1);
        _maxi_wstrb_sb_0 <= { 4{ 1'd1 } };
      end 
      _maxi_wdata_cond_1_1 <= 1;
      if(_maxi_wvalid_sb_0 && !_maxi_wready_sb_0) begin
        _maxi_wvalid_sb_0 <= _maxi_wvalid_sb_0;
        _maxi_wlast_sb_0 <= _maxi_wlast_sb_0;
      end 
      if((_maxi_write_op_sel_buf == 3) && read_burst_rvalid_1199 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0)) begin
        _maxi_wdata_sb_0 <= read_burst_rdata_1203;
        _maxi_wvalid_sb_0 <= 1;
        _maxi_wlast_sb_0 <= read_burst_rlast_1200 || (_maxi_write_size_buf == 1);
        _maxi_wstrb_sb_0 <= { 4{ 1'd1 } };
      end 
      _maxi_wdata_cond_2_1 <= 1;
      if(_maxi_wvalid_sb_0 && !_maxi_wready_sb_0) begin
        _maxi_wvalid_sb_0 <= _maxi_wvalid_sb_0;
        _maxi_wlast_sb_0 <= _maxi_wlast_sb_0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _sb_maxi_writedata_data_6 <= 0;
      _sb_maxi_writedata_valid_7 <= 0;
      _sb_maxi_writedata_tmp_data_9 <= 0;
      _sb_maxi_writedata_tmp_valid_10 <= 0;
    end else begin
      if(_sb_maxi_writedata_m_ready_5 || !_sb_maxi_writedata_valid_7) begin
        _sb_maxi_writedata_data_6 <= _sb_maxi_writedata_next_data_11;
        _sb_maxi_writedata_valid_7 <= _sb_maxi_writedata_next_valid_12;
      end 
      if(!_sb_maxi_writedata_tmp_valid_10 && _sb_maxi_writedata_valid_7 && !_sb_maxi_writedata_m_ready_5) begin
        _sb_maxi_writedata_tmp_data_9 <= _sb_maxi_writedata_s_data_3;
        _sb_maxi_writedata_tmp_valid_10 <= _sb_maxi_writedata_s_valid_4;
      end 
      if(_sb_maxi_writedata_tmp_valid_10 && _sb_maxi_writedata_m_ready_5) begin
        _sb_maxi_writedata_tmp_valid_10 <= 0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      maxi_araddr <= 0;
      maxi_arlen <= 0;
      maxi_arvalid <= 0;
      _maxi_raddr_cond_0_1 <= 0;
    end else begin
      if(_maxi_raddr_cond_0_1) begin
        maxi_arvalid <= 0;
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid)) begin
        maxi_araddr <= _maxi_read_global_addr;
        maxi_arlen <= _maxi_read_cur_global_size - 1;
        maxi_arvalid <= 1;
      end 
      _maxi_raddr_cond_0_1 <= 1;
      if(maxi_arvalid && !maxi_arready) begin
        maxi_arvalid <= maxi_arvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _sb_maxi_readdata_data_21 <= 0;
      _sb_maxi_readdata_valid_22 <= 0;
      _sb_maxi_readdata_tmp_data_24 <= 0;
      _sb_maxi_readdata_tmp_valid_25 <= 0;
    end else begin
      if(_sb_maxi_readdata_m_ready_20 || !_sb_maxi_readdata_valid_22) begin
        _sb_maxi_readdata_data_21 <= _sb_maxi_readdata_next_data_26;
        _sb_maxi_readdata_valid_22 <= _sb_maxi_readdata_next_valid_27;
      end 
      if(!_sb_maxi_readdata_tmp_valid_25 && _sb_maxi_readdata_valid_22 && !_sb_maxi_readdata_m_ready_20) begin
        _sb_maxi_readdata_tmp_data_24 <= _sb_maxi_readdata_s_data_18;
        _sb_maxi_readdata_tmp_valid_25 <= _sb_maxi_readdata_s_valid_19;
      end 
      if(_sb_maxi_readdata_tmp_valid_25 && _sb_maxi_readdata_m_ready_20) begin
        _sb_maxi_readdata_tmp_valid_25 <= 0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_outstanding_wcount <= 0;
      _maxi_read_start <= 0;
      _maxi_write_start <= 0;
      _maxi_global_base_addr <= 0;
      _maxi_read_op_sel <= 0;
      _maxi_read_global_addr <= 0;
      _maxi_read_global_size <= 0;
      _maxi_read_local_addr <= 0;
      _maxi_read_local_stride <= 0;
      _maxi_read_local_size <= 0;
      _maxi_read_local_blocksize <= 0;
      _maxi_read_req_busy <= 0;
      _maxi_read_cur_global_size <= 0;
      _maxi_read_data_busy <= 0;
      _maxi_read_op_sel_buf <= 0;
      _maxi_read_local_addr_buf <= 0;
      _maxi_read_local_stride_buf <= 0;
      _maxi_read_local_size_buf <= 0;
      _maxi_read_local_blocksize_buf <= 0;
      _maxi_write_op_sel <= 0;
      _maxi_write_global_addr <= 0;
      _maxi_write_global_size <= 0;
      _maxi_write_local_addr <= 0;
      _maxi_write_local_stride <= 0;
      _maxi_write_local_size <= 0;
      _maxi_write_local_blocksize <= 0;
      _maxi_write_req_busy <= 0;
      _maxi_write_cur_global_size <= 0;
      _maxi_write_data_busy <= 0;
      _maxi_write_op_sel_buf <= 0;
      _maxi_write_local_addr_buf <= 0;
      _maxi_write_local_stride_buf <= 0;
      _maxi_write_size_buf <= 0;
      _maxi_write_local_blocksize_buf <= 0;
    end else begin
      if(maxi_awvalid && maxi_awready && !(maxi_bvalid && maxi_bready) && (_maxi_outstanding_wcount < 7)) begin
        _maxi_outstanding_wcount <= _maxi_outstanding_wcount + 1;
      end 
      if(!(maxi_awvalid && maxi_awready) && (maxi_bvalid && maxi_bready) && (_maxi_outstanding_wcount > 0)) begin
        _maxi_outstanding_wcount <= _maxi_outstanding_wcount - 1;
      end 
      _maxi_read_start <= 0;
      _maxi_write_start <= 0;
      _maxi_global_base_addr <= _saxi_register_32;
      if((control_conv2d_25 == 2) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 1;
        _maxi_read_global_addr <= mask_addr_masked_55;
        _maxi_read_global_size <= cparam_conv2d_25_bias_num;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_conv2d_25_bias_num;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_req_fsm == 0) && _maxi_read_start) begin
        _maxi_read_req_busy <= 1;
      end 
      if(_maxi_read_start && _maxi_read_req_fifo_almost_full) begin
        _maxi_read_start <= 1;
      end 
      if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && (_maxi_read_global_size <= 256) && ((mask_addr_masked_65 & 4095) + (_maxi_read_global_size << 2) >= 4096)) begin
        _maxi_read_cur_global_size <= 4096 - (mask_addr_masked_67 & 4095) >> 2;
        _maxi_read_global_size <= _maxi_read_global_size - (4096 - (mask_addr_masked_69 & 4095) >> 2);
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && (_maxi_read_global_size <= 256)) begin
        _maxi_read_cur_global_size <= _maxi_read_global_size;
        _maxi_read_global_size <= 0;
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && ((mask_addr_masked_71 & 4095) + 1024 >= 4096)) begin
        _maxi_read_cur_global_size <= 4096 - (mask_addr_masked_73 & 4095) >> 2;
        _maxi_read_global_size <= _maxi_read_global_size - (4096 - (mask_addr_masked_75 & 4095) >> 2);
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full) begin
        _maxi_read_cur_global_size <= 256;
        _maxi_read_global_size <= _maxi_read_global_size - 256;
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid)) begin
        _maxi_read_global_addr <= _maxi_read_global_addr + (_maxi_read_cur_global_size << 2);
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid) && (_maxi_read_global_size == 0)) begin
        _maxi_read_req_busy <= 0;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_25 == 4) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 2;
        _maxi_read_global_addr <= mask_addr_masked_81;
        _maxi_read_global_size <= cparam_conv2d_25_scale_num;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_conv2d_25_scale_num;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_25 == 8) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 3;
        _maxi_read_global_addr <= mask_addr_masked_87;
        _maxi_read_global_size <= cparam_conv2d_25_filter_read_size;
        _maxi_read_local_addr <= conv2d_25_filter_page_dma_offset;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_conv2d_25_filter_read_size;
        _maxi_read_local_blocksize <= cparam_conv2d_25_filter_read_block;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_25 == 14) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 4;
        _maxi_read_global_addr <= mask_addr_masked_147;
        _maxi_read_global_size <= cparam_conv2d_25_act_read_size;
        _maxi_read_local_addr <= conv2d_25_act_page_dma_offset_0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_conv2d_25_act_read_size;
        _maxi_read_local_blocksize <= cparam_conv2d_25_act_read_block;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_25 == 17) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 5;
        _maxi_read_global_addr <= mask_addr_masked_171;
        _maxi_read_global_size <= cparam_conv2d_25_act_read_size;
        _maxi_read_local_addr <= conv2d_25_act_page_dma_offset_1;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_conv2d_25_act_read_size;
        _maxi_read_local_blocksize <= cparam_conv2d_25_act_read_block;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_25 == 20) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 6;
        _maxi_read_global_addr <= mask_addr_masked_195;
        _maxi_read_global_size <= cparam_conv2d_25_act_read_size;
        _maxi_read_local_addr <= conv2d_25_act_page_dma_offset_2;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_conv2d_25_act_read_size;
        _maxi_read_local_blocksize <= cparam_conv2d_25_act_read_block;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 6))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_25 == 29) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 1;
        _maxi_write_global_addr <= mask_addr_masked_921;
        _maxi_write_global_size <= conv2d_25_next_out_write_size;
        _maxi_write_local_addr <= conv2d_25_out_laddr_offset + conv2d_25_out_page_dma_offset;
        _maxi_write_local_stride <= 1;
        _maxi_write_local_size <= conv2d_25_next_out_write_size;
        _maxi_write_local_blocksize <= 1;
      end 
      if((_maxi_write_req_fsm == 0) && _maxi_write_start) begin
        _maxi_write_req_busy <= 1;
      end 
      if(_maxi_write_start && _maxi_write_req_fifo_almost_full) begin
        _maxi_write_start <= 1;
      end 
      if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && (_maxi_write_global_size <= 256) && ((mask_addr_masked_931 & 4095) + (_maxi_write_global_size << 2) >= 4096)) begin
        _maxi_write_cur_global_size <= 4096 - (mask_addr_masked_933 & 4095) >> 2;
        _maxi_write_global_size <= _maxi_write_global_size - (4096 - (mask_addr_masked_935 & 4095) >> 2);
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && (_maxi_write_global_size <= 256)) begin
        _maxi_write_cur_global_size <= _maxi_write_global_size;
        _maxi_write_global_size <= 0;
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && ((mask_addr_masked_937 & 4095) + 1024 >= 4096)) begin
        _maxi_write_cur_global_size <= 4096 - (mask_addr_masked_939 & 4095) >> 2;
        _maxi_write_global_size <= _maxi_write_global_size - (4096 - (mask_addr_masked_941 & 4095) >> 2);
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full) begin
        _maxi_write_cur_global_size <= 256;
        _maxi_write_global_size <= _maxi_write_global_size - 256;
      end 
      if((_maxi_write_req_fsm == 1) && ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6))) begin
        _maxi_write_global_addr <= _maxi_write_global_addr + (_maxi_write_cur_global_size << 2);
      end 
      if((_maxi_write_req_fsm == 1) && ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6)) && (_maxi_write_global_size == 0)) begin
        _maxi_write_req_busy <= 0;
      end 
      if((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1))) begin
        _maxi_write_data_busy <= 1;
        _maxi_write_op_sel_buf <= _maxi_write_op_sel_fifo;
        _maxi_write_local_addr_buf <= _maxi_write_local_addr_fifo;
        _maxi_write_local_stride_buf <= _maxi_write_local_stride_fifo;
        _maxi_write_size_buf <= _maxi_write_size_fifo;
        _maxi_write_local_blocksize_buf <= _maxi_write_local_blocksize_fifo;
      end 
      if(_maxi_write_data_fsm == 1) begin
        _maxi_write_size_buf <= 0;
      end 
      if((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_fifo;
      end 
      if((_maxi_write_data_fsm == 2) && read_burst_rvalid_953 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_buf - 1;
      end 
      if((_maxi_write_data_fsm == 2) && ((_maxi_write_op_sel_buf == 1) && read_burst_rvalid_953 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) && read_burst_rlast_954) begin
        _maxi_write_data_busy <= 0;
      end 
      if((control_max_pool_serial_27 == 5) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 7;
        _maxi_read_global_addr <= mask_addr_masked_959;
        _maxi_read_global_size <= cparam_max_pool_serial_27_act_read_size;
        _maxi_read_local_addr <= max_pool_serial_27_act_page_dma_offset;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_max_pool_serial_27_act_read_size;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 7))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_max_pool_serial_27 == 8) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 7;
        _maxi_read_global_addr <= mask_addr_masked_965;
        _maxi_read_global_size <= cparam_max_pool_serial_27_act_read_size;
        _maxi_read_local_addr <= max_pool_serial_27_act_page_dma_offset + cparam_max_pool_serial_27_act_read_size;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_max_pool_serial_27_act_read_size;
        _maxi_read_local_blocksize <= 1;
      end 
      if((control_max_pool_serial_27 == 15) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 2;
        _maxi_write_global_addr <= mask_addr_masked_1055;
        _maxi_write_global_size <= cparam_max_pool_serial_27_out_write_size;
        _maxi_write_local_addr <= max_pool_serial_27_out_page_dma_offset;
        _maxi_write_local_stride <= 1;
        _maxi_write_local_size <= cparam_max_pool_serial_27_out_write_size;
        _maxi_write_local_blocksize <= 1;
      end 
      if((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2))) begin
        _maxi_write_data_busy <= 1;
        _maxi_write_op_sel_buf <= _maxi_write_op_sel_fifo;
        _maxi_write_local_addr_buf <= _maxi_write_local_addr_fifo;
        _maxi_write_local_stride_buf <= _maxi_write_local_stride_fifo;
        _maxi_write_size_buf <= _maxi_write_size_fifo;
        _maxi_write_local_blocksize_buf <= _maxi_write_local_blocksize_fifo;
      end 
      if(_maxi_write_data_fsm == 1) begin
        _maxi_write_size_buf <= 0;
      end 
      if((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_fifo;
      end 
      if((_maxi_write_data_fsm == 2) && read_burst_rvalid_1059 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_buf - 1;
      end 
      if((_maxi_write_data_fsm == 2) && ((_maxi_write_op_sel_buf == 2) && read_burst_rvalid_1059 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) && read_burst_rlast_1060) begin
        _maxi_write_data_busy <= 0;
      end 
      if((control_max_pool_47 == 5) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 8;
        _maxi_read_global_addr <= mask_addr_masked_1065;
        _maxi_read_global_size <= cparam_max_pool_47_act_read_size;
        _maxi_read_local_addr <= max_pool_47_act_page_dma_offset_0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_max_pool_47_act_read_size;
        _maxi_read_local_blocksize <= cparam_max_pool_47_act_read_block;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 8))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_max_pool_47 == 8) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 9;
        _maxi_read_global_addr <= mask_addr_masked_1083;
        _maxi_read_global_size <= cparam_max_pool_47_act_read_size;
        _maxi_read_local_addr <= max_pool_47_act_page_dma_offset_1;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_max_pool_47_act_read_size;
        _maxi_read_local_blocksize <= cparam_max_pool_47_act_read_block;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 9))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_max_pool_47 == 15) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 3;
        _maxi_write_global_addr <= mask_addr_masked_1195;
        _maxi_write_global_size <= cparam_max_pool_47_out_write_size;
        _maxi_write_local_addr <= max_pool_47_out_page_dma_offset;
        _maxi_write_local_stride <= 1;
        _maxi_write_local_size <= cparam_max_pool_47_out_write_size;
        _maxi_write_local_blocksize <= 1;
      end 
      if((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 3))) begin
        _maxi_write_data_busy <= 1;
        _maxi_write_op_sel_buf <= _maxi_write_op_sel_fifo;
        _maxi_write_local_addr_buf <= _maxi_write_local_addr_fifo;
        _maxi_write_local_stride_buf <= _maxi_write_local_stride_fifo;
        _maxi_write_size_buf <= _maxi_write_size_fifo;
        _maxi_write_local_blocksize_buf <= _maxi_write_local_blocksize_fifo;
      end 
      if(_maxi_write_data_fsm == 1) begin
        _maxi_write_size_buf <= 0;
      end 
      if((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_fifo;
      end 
      if((_maxi_write_data_fsm == 2) && read_burst_rvalid_1199 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_buf - 1;
      end 
      if((_maxi_write_data_fsm == 2) && ((_maxi_write_op_sel_buf == 3) && read_burst_rvalid_1199 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) && read_burst_rlast_1200) begin
        _maxi_write_data_busy <= 0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      count__maxi_read_req_fifo <= 0;
      __tmp_63_1 <= 0;
    end else begin
      if(_maxi_read_req_fifo_enq && !_maxi_read_req_fifo_full && (_maxi_read_req_fifo_deq && !_maxi_read_req_fifo_empty)) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo;
      end else if(_maxi_read_req_fifo_enq && !_maxi_read_req_fifo_full) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo + 1;
      end else if(_maxi_read_req_fifo_deq && !_maxi_read_req_fifo_empty) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo - 1;
      end 
      __tmp_63_1 <= _tmp_63;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      count__maxi_write_req_fifo <= 0;
      __tmp_929_1 <= 0;
      __tmp_949_1 <= 0;
    end else begin
      if(_maxi_write_req_fifo_enq && !_maxi_write_req_fifo_full && (_maxi_write_req_fifo_deq && !_maxi_write_req_fifo_empty)) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo;
      end else if(_maxi_write_req_fifo_enq && !_maxi_write_req_fifo_full) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo + 1;
      end else if(_maxi_write_req_fifo_deq && !_maxi_write_req_fifo_empty) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo - 1;
      end 
      __tmp_929_1 <= _tmp_929;
      __tmp_949_1 <= _tmp_949;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      saxi_rdata <= 0;
      saxi_rvalid <= 0;
      _saxi_rdata_cond_0_1 <= 0;
    end else begin
      if(_saxi_rdata_cond_0_1) begin
        saxi_rvalid <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid)) begin
        saxi_rdata <= axislite_rdata_46;
        saxi_rvalid <= 1;
      end 
      _saxi_rdata_cond_0_1 <= 1;
      if(saxi_rvalid && !saxi_rready) begin
        saxi_rvalid <= saxi_rvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      saxi_bvalid <= 0;
      prev_awvalid_43 <= 0;
      prev_arvalid_44 <= 0;
      writevalid_41 <= 0;
      readvalid_42 <= 0;
      addr_40 <= 0;
      _saxi_register_0 <= 0;
      _saxi_flag_0 <= 0;
      _saxi_register_1 <= 0;
      _saxi_flag_1 <= 0;
      _saxi_register_2 <= 0;
      _saxi_flag_2 <= 0;
      _saxi_register_3 <= 0;
      _saxi_flag_3 <= 0;
      _saxi_register_4 <= 0;
      _saxi_flag_4 <= 0;
      _saxi_register_5 <= 0;
      _saxi_flag_5 <= 0;
      _saxi_register_6 <= 0;
      _saxi_flag_6 <= 0;
      _saxi_register_7 <= 0;
      _saxi_flag_7 <= 0;
      _saxi_register_8 <= 0;
      _saxi_flag_8 <= 0;
      _saxi_register_9 <= 0;
      _saxi_flag_9 <= 0;
      _saxi_register_10 <= 0;
      _saxi_flag_10 <= 0;
      _saxi_register_11 <= 0;
      _saxi_flag_11 <= 0;
      _saxi_register_12 <= 0;
      _saxi_flag_12 <= 0;
      _saxi_register_13 <= 0;
      _saxi_flag_13 <= 0;
      _saxi_register_14 <= 0;
      _saxi_flag_14 <= 0;
      _saxi_register_15 <= 0;
      _saxi_flag_15 <= 0;
      _saxi_register_16 <= 0;
      _saxi_flag_16 <= 0;
      _saxi_register_17 <= 0;
      _saxi_flag_17 <= 0;
      _saxi_register_18 <= 0;
      _saxi_flag_18 <= 0;
      _saxi_register_19 <= 0;
      _saxi_flag_19 <= 0;
      _saxi_register_20 <= 0;
      _saxi_flag_20 <= 0;
      _saxi_register_21 <= 0;
      _saxi_flag_21 <= 0;
      _saxi_register_22 <= 0;
      _saxi_flag_22 <= 0;
      _saxi_register_23 <= 0;
      _saxi_flag_23 <= 0;
      _saxi_register_24 <= 0;
      _saxi_flag_24 <= 0;
      _saxi_register_25 <= 0;
      _saxi_flag_25 <= 0;
      _saxi_register_26 <= 0;
      _saxi_flag_26 <= 0;
      _saxi_register_27 <= 0;
      _saxi_flag_27 <= 0;
      _saxi_register_28 <= 0;
      _saxi_flag_28 <= 0;
      _saxi_register_29 <= 0;
      _saxi_flag_29 <= 0;
      _saxi_register_30 <= 0;
      _saxi_flag_30 <= 0;
      _saxi_register_31 <= 55301184;
      _saxi_flag_31 <= 0;
      _saxi_register_32 <= 0;
      _saxi_flag_32 <= 0;
      _saxi_register_33 <= 27836480;
      _saxi_flag_33 <= 0;
      _saxi_register_34 <= 0;
      _saxi_flag_34 <= 0;
      _saxi_register_35 <= 589824;
      _saxi_flag_35 <= 0;
      _saxi_register_36 <= 2666496;
      _saxi_flag_36 <= 0;
      _saxi_register_11[0] <= (0 >> 0) & 1'd1;
      _saxi_register_9[0] <= (0 >> 0) & 1'd1;
      _saxi_register_11[1] <= (0 >> 1) & 1'd1;
      _saxi_register_9[1] <= (0 >> 1) & 1'd1;
      _saxi_register_11[2] <= (0 >> 2) & 1'd1;
      _saxi_register_9[2] <= (0 >> 2) & 1'd1;
      _saxi_register_11[3] <= (0 >> 3) & 1'd1;
      _saxi_register_9[3] <= (0 >> 3) & 1'd1;
      _saxi_register_11[4] <= (0 >> 4) & 1'd1;
      _saxi_register_9[4] <= (0 >> 4) & 1'd1;
      _saxi_register_11[5] <= (0 >> 5) & 1'd1;
      _saxi_register_9[5] <= (0 >> 5) & 1'd1;
      _saxi_register_11[6] <= (0 >> 6) & 1'd1;
      _saxi_register_9[6] <= (0 >> 6) & 1'd1;
      _saxi_register_11[7] <= (0 >> 7) & 1'd1;
      _saxi_register_9[7] <= (0 >> 7) & 1'd1;
      _saxi_register_11[8] <= (0 >> 8) & 1'd1;
      _saxi_register_9[8] <= (0 >> 8) & 1'd1;
      _saxi_register_11[9] <= (0 >> 9) & 1'd1;
      _saxi_register_9[9] <= (0 >> 9) & 1'd1;
      _saxi_register_11[10] <= (0 >> 10) & 1'd1;
      _saxi_register_9[10] <= (0 >> 10) & 1'd1;
      _saxi_register_11[11] <= (0 >> 11) & 1'd1;
      _saxi_register_9[11] <= (0 >> 11) & 1'd1;
      _saxi_register_11[12] <= (0 >> 12) & 1'd1;
      _saxi_register_9[12] <= (0 >> 12) & 1'd1;
      _saxi_register_11[13] <= (0 >> 13) & 1'd1;
      _saxi_register_9[13] <= (0 >> 13) & 1'd1;
      _saxi_register_11[14] <= (0 >> 14) & 1'd1;
      _saxi_register_9[14] <= (0 >> 14) & 1'd1;
      _saxi_register_11[15] <= (0 >> 15) & 1'd1;
      _saxi_register_9[15] <= (0 >> 15) & 1'd1;
      _saxi_register_11[16] <= (0 >> 16) & 1'd1;
      _saxi_register_9[16] <= (0 >> 16) & 1'd1;
      _saxi_register_11[17] <= (0 >> 17) & 1'd1;
      _saxi_register_9[17] <= (0 >> 17) & 1'd1;
      _saxi_register_11[18] <= (0 >> 18) & 1'd1;
      _saxi_register_9[18] <= (0 >> 18) & 1'd1;
      _saxi_register_11[19] <= (0 >> 19) & 1'd1;
      _saxi_register_9[19] <= (0 >> 19) & 1'd1;
      _saxi_register_11[20] <= (0 >> 20) & 1'd1;
      _saxi_register_9[20] <= (0 >> 20) & 1'd1;
      _saxi_register_11[21] <= (0 >> 21) & 1'd1;
      _saxi_register_9[21] <= (0 >> 21) & 1'd1;
      _saxi_register_11[22] <= (0 >> 22) & 1'd1;
      _saxi_register_9[22] <= (0 >> 22) & 1'd1;
      _saxi_register_11[23] <= (0 >> 23) & 1'd1;
      _saxi_register_9[23] <= (0 >> 23) & 1'd1;
      _saxi_register_11[24] <= (0 >> 24) & 1'd1;
      _saxi_register_9[24] <= (0 >> 24) & 1'd1;
      _saxi_register_11[25] <= (0 >> 25) & 1'd1;
      _saxi_register_9[25] <= (0 >> 25) & 1'd1;
      _saxi_register_11[26] <= (0 >> 26) & 1'd1;
      _saxi_register_9[26] <= (0 >> 26) & 1'd1;
      _saxi_register_11[27] <= (0 >> 27) & 1'd1;
      _saxi_register_9[27] <= (0 >> 27) & 1'd1;
      _saxi_register_11[28] <= (0 >> 28) & 1'd1;
      _saxi_register_9[28] <= (0 >> 28) & 1'd1;
      _saxi_register_11[29] <= (0 >> 29) & 1'd1;
      _saxi_register_9[29] <= (0 >> 29) & 1'd1;
      _saxi_register_11[30] <= (0 >> 30) & 1'd1;
      _saxi_register_9[30] <= (0 >> 30) & 1'd1;
      _saxi_register_11[31] <= (0 >> 31) & 1'd1;
      _saxi_register_9[31] <= (0 >> 31) & 1'd1;
      internal_state_counter <= 0;
    end else begin
      if(saxi_bvalid && saxi_bready) begin
        saxi_bvalid <= 0;
      end 
      if(saxi_wvalid && saxi_wready) begin
        saxi_bvalid <= 1;
      end 
      prev_awvalid_43 <= saxi_awvalid;
      prev_arvalid_44 <= saxi_arvalid;
      writevalid_41 <= 0;
      readvalid_42 <= 0;
      if(saxi_awready && saxi_awvalid && !saxi_bvalid) begin
        addr_40 <= saxi_awaddr;
        writevalid_41 <= 1;
      end else if(saxi_arready && saxi_arvalid) begin
        addr_40 <= saxi_araddr;
        readvalid_42 <= 1;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 0)) begin
        _saxi_register_0 <= axislite_resetval_48;
        _saxi_flag_0 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 1)) begin
        _saxi_register_1 <= axislite_resetval_48;
        _saxi_flag_1 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 2)) begin
        _saxi_register_2 <= axislite_resetval_48;
        _saxi_flag_2 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 3)) begin
        _saxi_register_3 <= axislite_resetval_48;
        _saxi_flag_3 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 4)) begin
        _saxi_register_4 <= axislite_resetval_48;
        _saxi_flag_4 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 5)) begin
        _saxi_register_5 <= axislite_resetval_48;
        _saxi_flag_5 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 6)) begin
        _saxi_register_6 <= axislite_resetval_48;
        _saxi_flag_6 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 7)) begin
        _saxi_register_7 <= axislite_resetval_48;
        _saxi_flag_7 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 8)) begin
        _saxi_register_8 <= axislite_resetval_48;
        _saxi_flag_8 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 9)) begin
        _saxi_register_9 <= axislite_resetval_48;
        _saxi_flag_9 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 10)) begin
        _saxi_register_10 <= axislite_resetval_48;
        _saxi_flag_10 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 11)) begin
        _saxi_register_11 <= axislite_resetval_48;
        _saxi_flag_11 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 12)) begin
        _saxi_register_12 <= axislite_resetval_48;
        _saxi_flag_12 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 13)) begin
        _saxi_register_13 <= axislite_resetval_48;
        _saxi_flag_13 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 14)) begin
        _saxi_register_14 <= axislite_resetval_48;
        _saxi_flag_14 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 15)) begin
        _saxi_register_15 <= axislite_resetval_48;
        _saxi_flag_15 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 16)) begin
        _saxi_register_16 <= axislite_resetval_48;
        _saxi_flag_16 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 17)) begin
        _saxi_register_17 <= axislite_resetval_48;
        _saxi_flag_17 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 18)) begin
        _saxi_register_18 <= axislite_resetval_48;
        _saxi_flag_18 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 19)) begin
        _saxi_register_19 <= axislite_resetval_48;
        _saxi_flag_19 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 20)) begin
        _saxi_register_20 <= axislite_resetval_48;
        _saxi_flag_20 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 21)) begin
        _saxi_register_21 <= axislite_resetval_48;
        _saxi_flag_21 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 22)) begin
        _saxi_register_22 <= axislite_resetval_48;
        _saxi_flag_22 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 23)) begin
        _saxi_register_23 <= axislite_resetval_48;
        _saxi_flag_23 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 24)) begin
        _saxi_register_24 <= axislite_resetval_48;
        _saxi_flag_24 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 25)) begin
        _saxi_register_25 <= axislite_resetval_48;
        _saxi_flag_25 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 26)) begin
        _saxi_register_26 <= axislite_resetval_48;
        _saxi_flag_26 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 27)) begin
        _saxi_register_27 <= axislite_resetval_48;
        _saxi_flag_27 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 28)) begin
        _saxi_register_28 <= axislite_resetval_48;
        _saxi_flag_28 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 29)) begin
        _saxi_register_29 <= axislite_resetval_48;
        _saxi_flag_29 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 30)) begin
        _saxi_register_30 <= axislite_resetval_48;
        _saxi_flag_30 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 31)) begin
        _saxi_register_31 <= axislite_resetval_48;
        _saxi_flag_31 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 32)) begin
        _saxi_register_32 <= axislite_resetval_48;
        _saxi_flag_32 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 33)) begin
        _saxi_register_33 <= axislite_resetval_48;
        _saxi_flag_33 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 34)) begin
        _saxi_register_34 <= axislite_resetval_48;
        _saxi_flag_34 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 35)) begin
        _saxi_register_35 <= axislite_resetval_48;
        _saxi_flag_35 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 36)) begin
        _saxi_register_36 <= axislite_resetval_48;
        _saxi_flag_36 <= 0;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 0)) begin
        _saxi_register_0 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 1)) begin
        _saxi_register_1 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 2)) begin
        _saxi_register_2 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 3)) begin
        _saxi_register_3 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 4)) begin
        _saxi_register_4 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 5)) begin
        _saxi_register_5 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 6)) begin
        _saxi_register_6 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 7)) begin
        _saxi_register_7 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 8)) begin
        _saxi_register_8 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 9)) begin
        _saxi_register_9 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 10)) begin
        _saxi_register_10 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 11)) begin
        _saxi_register_11 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 12)) begin
        _saxi_register_12 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 13)) begin
        _saxi_register_13 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 14)) begin
        _saxi_register_14 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 15)) begin
        _saxi_register_15 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 16)) begin
        _saxi_register_16 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 17)) begin
        _saxi_register_17 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 18)) begin
        _saxi_register_18 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 19)) begin
        _saxi_register_19 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 20)) begin
        _saxi_register_20 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 21)) begin
        _saxi_register_21 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 22)) begin
        _saxi_register_22 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 23)) begin
        _saxi_register_23 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 24)) begin
        _saxi_register_24 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 25)) begin
        _saxi_register_25 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 26)) begin
        _saxi_register_26 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 27)) begin
        _saxi_register_27 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 28)) begin
        _saxi_register_28 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 29)) begin
        _saxi_register_29 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 30)) begin
        _saxi_register_30 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 31)) begin
        _saxi_register_31 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 32)) begin
        _saxi_register_32 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 33)) begin
        _saxi_register_33 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 34)) begin
        _saxi_register_34 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 35)) begin
        _saxi_register_35 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 36)) begin
        _saxi_register_36 <= saxi_wdata;
      end 
      if(_saxi_register_11[0] == 1) begin
        _saxi_register_11[0] <= 0;
        _saxi_register_9[0] <= 0;
      end 
      if(_saxi_register_11[1] == 1) begin
        _saxi_register_11[1] <= 0;
        _saxi_register_9[1] <= 0;
      end 
      if(_saxi_register_11[2] == 1) begin
        _saxi_register_11[2] <= 0;
        _saxi_register_9[2] <= 0;
      end 
      if(_saxi_register_11[3] == 1) begin
        _saxi_register_11[3] <= 0;
        _saxi_register_9[3] <= 0;
      end 
      if(_saxi_register_11[4] == 1) begin
        _saxi_register_11[4] <= 0;
        _saxi_register_9[4] <= 0;
      end 
      if(_saxi_register_11[5] == 1) begin
        _saxi_register_11[5] <= 0;
        _saxi_register_9[5] <= 0;
      end 
      if(_saxi_register_11[6] == 1) begin
        _saxi_register_11[6] <= 0;
        _saxi_register_9[6] <= 0;
      end 
      if(_saxi_register_11[7] == 1) begin
        _saxi_register_11[7] <= 0;
        _saxi_register_9[7] <= 0;
      end 
      if(_saxi_register_11[8] == 1) begin
        _saxi_register_11[8] <= 0;
        _saxi_register_9[8] <= 0;
      end 
      if(_saxi_register_11[9] == 1) begin
        _saxi_register_11[9] <= 0;
        _saxi_register_9[9] <= 0;
      end 
      if(_saxi_register_11[10] == 1) begin
        _saxi_register_11[10] <= 0;
        _saxi_register_9[10] <= 0;
      end 
      if(_saxi_register_11[11] == 1) begin
        _saxi_register_11[11] <= 0;
        _saxi_register_9[11] <= 0;
      end 
      if(_saxi_register_11[12] == 1) begin
        _saxi_register_11[12] <= 0;
        _saxi_register_9[12] <= 0;
      end 
      if(_saxi_register_11[13] == 1) begin
        _saxi_register_11[13] <= 0;
        _saxi_register_9[13] <= 0;
      end 
      if(_saxi_register_11[14] == 1) begin
        _saxi_register_11[14] <= 0;
        _saxi_register_9[14] <= 0;
      end 
      if(_saxi_register_11[15] == 1) begin
        _saxi_register_11[15] <= 0;
        _saxi_register_9[15] <= 0;
      end 
      if(_saxi_register_11[16] == 1) begin
        _saxi_register_11[16] <= 0;
        _saxi_register_9[16] <= 0;
      end 
      if(_saxi_register_11[17] == 1) begin
        _saxi_register_11[17] <= 0;
        _saxi_register_9[17] <= 0;
      end 
      if(_saxi_register_11[18] == 1) begin
        _saxi_register_11[18] <= 0;
        _saxi_register_9[18] <= 0;
      end 
      if(_saxi_register_11[19] == 1) begin
        _saxi_register_11[19] <= 0;
        _saxi_register_9[19] <= 0;
      end 
      if(_saxi_register_11[20] == 1) begin
        _saxi_register_11[20] <= 0;
        _saxi_register_9[20] <= 0;
      end 
      if(_saxi_register_11[21] == 1) begin
        _saxi_register_11[21] <= 0;
        _saxi_register_9[21] <= 0;
      end 
      if(_saxi_register_11[22] == 1) begin
        _saxi_register_11[22] <= 0;
        _saxi_register_9[22] <= 0;
      end 
      if(_saxi_register_11[23] == 1) begin
        _saxi_register_11[23] <= 0;
        _saxi_register_9[23] <= 0;
      end 
      if(_saxi_register_11[24] == 1) begin
        _saxi_register_11[24] <= 0;
        _saxi_register_9[24] <= 0;
      end 
      if(_saxi_register_11[25] == 1) begin
        _saxi_register_11[25] <= 0;
        _saxi_register_9[25] <= 0;
      end 
      if(_saxi_register_11[26] == 1) begin
        _saxi_register_11[26] <= 0;
        _saxi_register_9[26] <= 0;
      end 
      if(_saxi_register_11[27] == 1) begin
        _saxi_register_11[27] <= 0;
        _saxi_register_9[27] <= 0;
      end 
      if(_saxi_register_11[28] == 1) begin
        _saxi_register_11[28] <= 0;
        _saxi_register_9[28] <= 0;
      end 
      if(_saxi_register_11[29] == 1) begin
        _saxi_register_11[29] <= 0;
        _saxi_register_9[29] <= 0;
      end 
      if(_saxi_register_11[30] == 1) begin
        _saxi_register_11[30] <= 0;
        _saxi_register_9[30] <= 0;
      end 
      if(_saxi_register_11[31] == 1) begin
        _saxi_register_11[31] <= 0;
        _saxi_register_9[31] <= 0;
      end 
      if(irq_busy_edge_51) begin
        _saxi_register_9[0] <= irq_busy_edge_51;
      end 
      if(irq_extern_edge_53) begin
        _saxi_register_9[1] <= irq_extern_edge_53;
      end 
      if(main_fsm == 0) begin
        _saxi_register_5 <= 0;
        _saxi_register_6 <= 0;
        _saxi_register_7 <= 0;
      end 
      if(main_fsm == 1) begin
        internal_state_counter <= 0;
        _saxi_register_12 <= 0;
      end else if(main_fsm == _saxi_register_13) begin
        if(internal_state_counter == _saxi_register_14) begin
          internal_state_counter <= 0;
          _saxi_register_12 <= _saxi_register_12 + 1;
        end else begin
          internal_state_counter <= internal_state_counter + 1;
        end
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_0 <= 1;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_1 <= 1;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_2 <= 1;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_3 <= 1;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_4 <= 1;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 1) && 1) begin
        _saxi_register_5 <= 1;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_6 <= 1;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_7 <= 1;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_8 <= 1;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_9 <= 1;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_10 <= 1;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_11 <= 1;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_12 <= 1;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_13 <= 1;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_14 <= 1;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_15 <= 1;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_16 <= 1;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_17 <= 1;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_18 <= 1;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_19 <= 1;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_20 <= 1;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_21 <= 1;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_22 <= 1;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_23 <= 1;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_24 <= 1;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_25 <= 1;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_26 <= 1;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_27 <= 1;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_28 <= 1;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_29 <= 1;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_30 <= 1;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_31 <= 1;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_32 <= 1;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_33 <= 1;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_34 <= 1;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_35 <= 1;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_36 <= 1;
        _saxi_flag_36 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_0 <= 0;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_1 <= 0;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_2 <= 0;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_3 <= 0;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 2) && 1) begin
        _saxi_register_4 <= 0;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_5 <= 0;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_6 <= 0;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_7 <= 0;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_8 <= 0;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_9 <= 0;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_10 <= 0;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_11 <= 0;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_12 <= 0;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_13 <= 0;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_14 <= 0;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_15 <= 0;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_16 <= 0;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_17 <= 0;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_18 <= 0;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_19 <= 0;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_20 <= 0;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_21 <= 0;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_22 <= 0;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_23 <= 0;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_24 <= 0;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_25 <= 0;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_26 <= 0;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_27 <= 0;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_28 <= 0;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_29 <= 0;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_30 <= 0;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_31 <= 0;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_32 <= 0;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_33 <= 0;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_34 <= 0;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_35 <= 0;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_36 <= 0;
        _saxi_flag_36 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_0 <= 0;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_1 <= 0;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_2 <= 0;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_3 <= 0;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_4 <= 0;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 117) && 1) begin
        _saxi_register_5 <= 0;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_6 <= 0;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_7 <= 0;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_8 <= 0;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_9 <= 0;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_10 <= 0;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_11 <= 0;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_12 <= 0;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_13 <= 0;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_14 <= 0;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_15 <= 0;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_16 <= 0;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_17 <= 0;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_18 <= 0;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_19 <= 0;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_20 <= 0;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_21 <= 0;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_22 <= 0;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_23 <= 0;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_24 <= 0;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_25 <= 0;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_26 <= 0;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_27 <= 0;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_28 <= 0;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_29 <= 0;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_30 <= 0;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_31 <= 0;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_32 <= 0;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_33 <= 0;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_34 <= 0;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_35 <= 0;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 117) && 0) begin
        _saxi_register_36 <= 0;
        _saxi_flag_36 <= 0;
      end 
    end
  end

  localparam _saxi_register_fsm_1 = 1;
  localparam _saxi_register_fsm_2 = 2;
  localparam _saxi_register_fsm_3 = 3;
  localparam _saxi_register_fsm_4 = 4;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _saxi_register_fsm <= _saxi_register_fsm_init;
      axis_maskaddr_45 <= 0;
    end else begin
      case(_saxi_register_fsm)
        _saxi_register_fsm_init: begin
          if(readvalid_42 || writevalid_41) begin
            axis_maskaddr_45 <= (addr_40 >> _saxi_shift) & _saxi_mask;
          end 
          if(readvalid_42) begin
            _saxi_register_fsm <= _saxi_register_fsm_1;
          end 
          if(writevalid_41) begin
            _saxi_register_fsm <= _saxi_register_fsm_3;
          end 
        end
        _saxi_register_fsm_1: begin
          if(saxi_rready || !saxi_rvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_2;
          end 
        end
        _saxi_register_fsm_2: begin
          if(saxi_rready && saxi_rvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_init;
          end 
        end
        _saxi_register_fsm_3: begin
          if(saxi_wvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_4;
          end 
        end
        _saxi_register_fsm_4: begin
          if(saxi_bready && saxi_bvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    _rst_logic_1 <= rst_logic;
    _rst_logic_2 <= _rst_logic_1;
    RST <= rst_logic | _rst_logic_1 | _rst_logic_2;
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq <= 0;
    end else begin
      irq <= |irq_49;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq_busy_edge_50 <= 0;
    end else begin
      irq_busy_edge_50 <= irq_busy;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq_extern_edge_52 <= 0;
    end else begin
      irq_extern_edge_52 <= irq_extern;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_970_1 <= 0;
    end else begin
      __tmp_970_1 <= _tmp_970;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1202_1 <= 0;
    end else begin
      __tmp_1202_1 <= _tmp_1202;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_267_1 <= 0;
      __tmp_1062_1 <= 0;
      __tmp_1103_1 <= 0;
    end else begin
      __tmp_267_1 <= _tmp_267;
      __tmp_1062_1 <= _tmp_1062;
      __tmp_1103_1 <= _tmp_1103;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1106_1 <= 0;
    end else begin
      __tmp_1106_1 <= _tmp_1106;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1109_1 <= 0;
    end else begin
      __tmp_1109_1 <= _tmp_1109;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1112_1 <= 0;
    end else begin
      __tmp_1112_1 <= _tmp_1112;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_226_1 <= 0;
    end else begin
      __tmp_226_1 <= _tmp_226;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_243_1 <= 0;
    end else begin
      __tmp_243_1 <= _tmp_243;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_246_1 <= 0;
    end else begin
      __tmp_246_1 <= _tmp_246;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_249_1 <= 0;
    end else begin
      __tmp_249_1 <= _tmp_249;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_252_1 <= 0;
    end else begin
      __tmp_252_1 <= _tmp_252;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_255_1 <= 0;
    end else begin
      __tmp_255_1 <= _tmp_255;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_258_1 <= 0;
    end else begin
      __tmp_258_1 <= _tmp_258;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_261_1 <= 0;
    end else begin
      __tmp_261_1 <= _tmp_261;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_264_1 <= 0;
    end else begin
      __tmp_264_1 <= _tmp_264;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_230_1 <= 0;
    end else begin
      __tmp_230_1 <= _tmp_230;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_956_1 <= 0;
    end else begin
      __tmp_956_1 <= _tmp_956;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_270_1 <= 0;
    end else begin
      __tmp_270_1 <= _tmp_270;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_273_1 <= 0;
    end else begin
      __tmp_273_1 <= _tmp_273;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_276_1 <= 0;
    end else begin
      __tmp_276_1 <= _tmp_276;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_279_1 <= 0;
    end else begin
      __tmp_279_1 <= _tmp_279;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_282_1 <= 0;
    end else begin
      __tmp_282_1 <= _tmp_282;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_285_1 <= 0;
    end else begin
      __tmp_285_1 <= _tmp_285;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_288_1 <= 0;
    end else begin
      __tmp_288_1 <= _tmp_288;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_291_1 <= 0;
    end else begin
      __tmp_291_1 <= _tmp_291;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_294_1 <= 0;
    end else begin
      __tmp_294_1 <= _tmp_294;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __max_0_var0_source_ram_renable <= 0;
      __max_0_var0_source_fifo_deq <= 0;
      __max_0_var0_idle <= 1;
      __max_0_var1_source_ram_renable <= 0;
      __max_0_var1_source_fifo_deq <= 0;
      __max_0_var1_idle <= 1;
      __max_0_var2_source_ram_renable <= 0;
      __max_0_var2_source_fifo_deq <= 0;
      __max_0_var2_idle <= 1;
      __max_0_var3_source_ram_renable <= 0;
      __max_0_var3_source_fifo_deq <= 0;
      __max_0_var3_idle <= 1;
      __max_0_val_sink_wenable <= 0;
      __max_0_val_sink_fifo_enq <= 0;
      ___max_0_stream_ivalid_1 <= 0;
      ___max_0_stream_ivalid_2 <= 0;
      ___max_0_stream_ivalid_3 <= 0;
      ___max_0_stream_ivalid_4 <= 0;
      _greaterthan_data_4 <= 0;
      _greaterthan_data_6 <= 0;
      __delay_data_938__variable_0 <= 0;
      __delay_data_939__variable_1 <= 0;
      __delay_data_940__variable_2 <= 0;
      __delay_data_941__variable_3 <= 0;
      _cond_data_5 <= 0;
      _cond_data_7 <= 0;
      _greaterthan_data_8 <= 0;
      __delay_data_942_cond_5 <= 0;
      __delay_data_943_cond_7 <= 0;
      _cond_data_9 <= 0;
      __variable_wdata_0 <= 0;
      __variable_wdata_1 <= 0;
      __variable_wdata_2 <= 0;
      __variable_wdata_3 <= 0;
      _tmp_1141 <= 0;
      _tmp_1142 <= 0;
      _tmp_1143 <= 0;
      _tmp_1144 <= 0;
      _tmp_1145 <= 0;
      _tmp_1146 <= 0;
      _tmp_1147 <= 0;
      _tmp_1148 <= 0;
      _tmp_1149 <= 0;
      _tmp_1150 <= 0;
      _tmp_1151 <= 0;
      _tmp_1152 <= 0;
      _tmp_1153 <= 0;
      _tmp_1154 <= 0;
      _tmp_1155 <= 0;
      _tmp_1156 <= 0;
      _tmp_1157 <= 0;
      _tmp_1158 <= 0;
      _tmp_1159 <= 0;
      _tmp_1160 <= 0;
      _tmp_1161 <= 0;
      _tmp_1162 <= 0;
      __max_0_busy_reg <= 0;
    end else begin
      if(__max_0_stream_oready) begin
        __max_0_var0_source_ram_renable <= 0;
        __max_0_var0_source_fifo_deq <= 0;
      end 
      __max_0_var0_idle <= __max_0_var0_idle;
      if(__max_0_stream_oready) begin
        __max_0_var1_source_ram_renable <= 0;
        __max_0_var1_source_fifo_deq <= 0;
      end 
      __max_0_var1_idle <= __max_0_var1_idle;
      if(__max_0_stream_oready) begin
        __max_0_var2_source_ram_renable <= 0;
        __max_0_var2_source_fifo_deq <= 0;
      end 
      __max_0_var2_idle <= __max_0_var2_idle;
      if(__max_0_stream_oready) begin
        __max_0_var3_source_ram_renable <= 0;
        __max_0_var3_source_fifo_deq <= 0;
      end 
      __max_0_var3_idle <= __max_0_var3_idle;
      if(__max_0_stream_oready) begin
        __max_0_val_sink_wenable <= 0;
        __max_0_val_sink_fifo_enq <= 0;
      end 
      if(__max_0_stream_oready) begin
        ___max_0_stream_ivalid_1 <= __max_0_stream_ivalid;
      end 
      if(__max_0_stream_oready) begin
        ___max_0_stream_ivalid_2 <= ___max_0_stream_ivalid_1;
      end 
      if(__max_0_stream_oready) begin
        ___max_0_stream_ivalid_3 <= ___max_0_stream_ivalid_2;
      end 
      if(__max_0_stream_oready) begin
        ___max_0_stream_ivalid_4 <= ___max_0_stream_ivalid_3;
      end 
      if(__max_0_stream_oready) begin
        _greaterthan_data_4 <= _max_0_var0_data > _max_0_var1_data;
      end 
      if(__max_0_stream_oready) begin
        _greaterthan_data_6 <= _max_0_var2_data > _max_0_var3_data;
      end 
      if(__max_0_stream_oready) begin
        __delay_data_938__variable_0 <= _max_0_var0_data;
      end 
      if(__max_0_stream_oready) begin
        __delay_data_939__variable_1 <= _max_0_var1_data;
      end 
      if(__max_0_stream_oready) begin
        __delay_data_940__variable_2 <= _max_0_var2_data;
      end 
      if(__max_0_stream_oready) begin
        __delay_data_941__variable_3 <= _max_0_var3_data;
      end 
      if(__max_0_stream_oready) begin
        _cond_data_5 <= (_greaterthan_data_4)? __delay_data_938__variable_0 : __delay_data_939__variable_1;
      end 
      if(__max_0_stream_oready) begin
        _cond_data_7 <= (_greaterthan_data_6)? __delay_data_940__variable_2 : __delay_data_941__variable_3;
      end 
      if(__max_0_stream_oready) begin
        _greaterthan_data_8 <= _cond_data_5 > _cond_data_7;
      end 
      if(__max_0_stream_oready) begin
        __delay_data_942_cond_5 <= _cond_data_5;
      end 
      if(__max_0_stream_oready) begin
        __delay_data_943_cond_7 <= _cond_data_7;
      end 
      if(__max_0_stream_oready) begin
        _cond_data_9 <= (_greaterthan_data_8)? __delay_data_942_cond_5 : __delay_data_943_cond_7;
      end 
      if(__stream_max_pool_47_stream_ivalid_1 && _stream_max_pool_47_stream_oready) begin
        __variable_wdata_0 <= _cond_data_927;
      end 
      if(__stream_max_pool_47_stream_ivalid_1 && _stream_max_pool_47_stream_oready) begin
        __variable_wdata_1 <= _cond_data_930;
      end 
      if(__stream_max_pool_47_stream_ivalid_1 && _stream_max_pool_47_stream_oready) begin
        __variable_wdata_2 <= _cond_data_933;
      end 
      if(__stream_max_pool_47_stream_ivalid_1 && _stream_max_pool_47_stream_oready) begin
        __variable_wdata_3 <= _cond_data_936;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1141 <= __max_0_source_start;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1142 <= _tmp_1141;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1143 <= _tmp_1142;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1144 <= __max_0_source_start;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1145 <= _tmp_1144;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1146 <= _tmp_1145;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1147 <= _tmp_1146;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1148 <= _tmp_1147;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1149 <= _tmp_1148;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1150 <= __max_0_source_stop;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1151 <= _tmp_1150;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1152 <= _tmp_1151;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1153 <= _tmp_1152;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1154 <= _tmp_1153;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1155 <= _tmp_1154;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1156 <= __max_0_source_busy;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1157 <= _tmp_1156;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1158 <= _tmp_1157;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1159 <= _tmp_1158;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1160 <= _tmp_1159;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1161 <= _tmp_1160;
      end 
      if(__max_0_stream_oready) begin
        _tmp_1162 <= __max_0_sink_busy;
      end 
      if(!__max_0_sink_busy && _tmp_1162) begin
        __max_0_busy_reg <= 0;
      end 
      if(__max_0_source_busy) begin
        __max_0_busy_reg <= 1;
      end 
    end
  end

  localparam __max_0_fsm_1 = 1;
  localparam __max_0_fsm_2 = 2;
  localparam __max_0_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      __max_0_fsm <= __max_0_fsm_init;
      __max_0_source_start <= 0;
      __max_0_source_busy <= 0;
      __max_0_stream_ivalid <= 0;
    end else begin
      if(__stream_max_pool_47_stream_ivalid_1 && _stream_max_pool_47_stream_oready) begin
        __max_0_stream_ivalid <= 1'd1;
      end 
      if(_stream_max_pool_47_stream_oready && _stream_max_pool_47_busy) begin
        __max_0_source_busy <= _stream_max_pool_47_source_busy;
      end 
      if(__max_0_stream_oready && _tmp_1143) begin
        __max_0_stream_ivalid <= 1;
      end 
      if(__max_0_stream_oready && 1'd0) begin
        __max_0_stream_ivalid <= 0;
      end 
      case(__max_0_fsm)
        __max_0_fsm_init: begin
          if(__max_0_run_flag) begin
            __max_0_source_start <= 1;
          end 
          if(__max_0_run_flag) begin
            __max_0_fsm <= __max_0_fsm_1;
          end 
        end
        __max_0_fsm_1: begin
          if(__max_0_source_start && __max_0_stream_oready) begin
            __max_0_source_start <= 0;
            __max_0_source_busy <= 1;
          end 
          if(__max_0_source_start && __max_0_stream_oready) begin
            __max_0_fsm <= __max_0_fsm_2;
          end 
        end
        __max_0_fsm_2: begin
          if(__max_0_stream_oready) begin
            __max_0_fsm <= __max_0_fsm_3;
          end 
        end
        __max_0_fsm_3: begin
          if(__max_0_stream_oready && 1'd0) begin
            __max_0_source_busy <= 0;
          end 
          if(__max_0_stream_oready && 1'd0 && __max_0_run_flag) begin
            __max_0_source_start <= 1;
          end 
          if(__max_0_stream_oready && 1'd0) begin
            __max_0_fsm <= __max_0_fsm_init;
          end 
          if(__max_0_stream_oready && 1'd0 && __max_0_run_flag) begin
            __max_0_fsm <= __max_0_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _acc_1_x_source_ram_renable <= 0;
      _acc_1_x_source_fifo_deq <= 0;
      _acc_1_x_idle <= 1;
      _acc_1_rshift_source_ram_renable <= 0;
      _acc_1_rshift_source_fifo_deq <= 0;
      _acc_1_rshift_idle <= 1;
      _acc_1_sum_sink_wenable <= 0;
      _acc_1_sum_sink_fifo_enq <= 0;
      _acc_1_valid_sink_wenable <= 0;
      _acc_1_valid_sink_fifo_enq <= 0;
      __acc_1_stream_ivalid_1 <= 0;
      __acc_1_stream_ivalid_2 <= 0;
      __acc_1_stream_ivalid_3 <= 0;
      __acc_1_stream_ivalid_4 <= 0;
      __acc_1_stream_ivalid_5 <= 0;
      _greaterthan_data_13 <= 0;
      _minus_data_15 <= 0;
      _reduceadd_data_26 <= 1'sd0;
      _reduceadd_count_26 <= 0;
      _reduceadd_prev_count_max_26 <= 0;
      _pulse_data_28 <= 1'sd0;
      _pulse_count_28 <= 0;
      _pulse_prev_count_max_28 <= 0;
      __delay_data_831__variable_11 <= 0;
      _sll_data_17 <= 0;
      __delay_data_828_greaterthan_13 <= 0;
      __delay_data_829_reduceadd_26 <= 0;
      __delay_data_832__delay_831__variable_11 <= 0;
      __delay_data_835_pulse_28 <= 0;
      _cond_data_23 <= 0;
      __delay_data_830__delay_829_reduceadd_26 <= 0;
      __delay_data_833__delay_832__delay_831__variable_11 <= 0;
      __delay_data_836__delay_835_pulse_28 <= 0;
      _plus_data_30 <= 0;
      __delay_data_834__delay_833__delay_832__delay_831__variable_11 <= 0;
      __delay_data_837__delay_836__delay_835_pulse_28 <= 0;
      _sra_data_31 <= 0;
      __delay_data_838__delay_837__delay_836__delay_835_pulse_28 <= 0;
      __variable_wdata_25 <= 0;
      __variable_wdata_10 <= 0;
      __variable_wdata_11 <= 0;
      __variable_wdata_12 <= 0;
      _tmp_729 <= 0;
      _tmp_730 <= 0;
      _tmp_731 <= 0;
      _tmp_732 <= 0;
      _tmp_733 <= 0;
      _tmp_734 <= 0;
      _tmp_735 <= 0;
      _tmp_736 <= 0;
      _tmp_737 <= 0;
      _tmp_738 <= 0;
      _tmp_739 <= 0;
      _tmp_740 <= 0;
      _tmp_741 <= 0;
      _tmp_742 <= 0;
      _tmp_743 <= 0;
      _tmp_744 <= 0;
      _tmp_745 <= 0;
      _tmp_746 <= 0;
      _tmp_747 <= 0;
      _tmp_748 <= 0;
      _tmp_749 <= 0;
      _tmp_750 <= 0;
      _tmp_751 <= 0;
      _tmp_752 <= 0;
      _tmp_753 <= 0;
      _tmp_754 <= 0;
      _tmp_755 <= 0;
      _tmp_756 <= 0;
      _tmp_757 <= 0;
      _tmp_758 <= 0;
      _tmp_759 <= 0;
      _tmp_760 <= 0;
      _acc_1_busy_reg <= 0;
    end else begin
      if(_acc_1_stream_oready) begin
        _acc_1_x_source_ram_renable <= 0;
        _acc_1_x_source_fifo_deq <= 0;
      end 
      _acc_1_x_idle <= _acc_1_x_idle;
      if(_acc_1_stream_oready) begin
        _acc_1_rshift_source_ram_renable <= 0;
        _acc_1_rshift_source_fifo_deq <= 0;
      end 
      _acc_1_rshift_idle <= _acc_1_rshift_idle;
      if(_acc_1_stream_oready) begin
        _acc_1_sum_sink_wenable <= 0;
        _acc_1_sum_sink_fifo_enq <= 0;
      end 
      if(_acc_1_stream_oready) begin
        _acc_1_valid_sink_wenable <= 0;
        _acc_1_valid_sink_fifo_enq <= 0;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_1 <= _acc_1_stream_ivalid;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_2 <= __acc_1_stream_ivalid_1;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_3 <= __acc_1_stream_ivalid_2;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_4 <= __acc_1_stream_ivalid_3;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_5 <= __acc_1_stream_ivalid_4;
      end 
      if(_acc_1_stream_oready) begin
        _greaterthan_data_13 <= acc_1_rshift_data > 1'sd0;
      end 
      if(_acc_1_stream_oready) begin
        _minus_data_15 <= acc_1_rshift_data - 2'sd1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready && _reduceadd_reset_cond_26) begin
        _reduceadd_data_26 <= 1'sd0;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _reduceadd_count_26 <= (_reduceadd_current_count_26 >= acc_1_size_data - 1)? 0 : _reduceadd_current_count_26 + 1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _reduceadd_prev_count_max_26 <= _reduceadd_current_count_26 >= acc_1_size_data - 1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _reduceadd_data_26 <= _reduceadd_current_data_26 + acc_1_x_data;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready && _pulse_reset_cond_28) begin
        _pulse_data_28 <= 1'sd0;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _pulse_count_28 <= (_pulse_current_count_28 >= acc_1_size_data - 1)? 0 : _pulse_current_count_28 + 1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _pulse_prev_count_max_28 <= _pulse_current_count_28 >= acc_1_size_data - 1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _pulse_data_28 <= _pulse_current_count_28 >= acc_1_size_data - 1;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_831__variable_11 <= acc_1_rshift_data;
      end 
      if(_acc_1_stream_oready) begin
        _sll_data_17 <= 2'sd1 << _minus_data_15;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_828_greaterthan_13 <= _greaterthan_data_13;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_829_reduceadd_26 <= _reduceadd_data_26;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_832__delay_831__variable_11 <= __delay_data_831__variable_11;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_835_pulse_28 <= _pulse_data_28;
      end 
      if(_acc_1_stream_oready) begin
        _cond_data_23 <= (__delay_data_828_greaterthan_13)? _sll_data_17 : 1'sd0;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_830__delay_829_reduceadd_26 <= __delay_data_829_reduceadd_26;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_833__delay_832__delay_831__variable_11 <= __delay_data_832__delay_831__variable_11;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_836__delay_835_pulse_28 <= __delay_data_835_pulse_28;
      end 
      if(_acc_1_stream_oready) begin
        _plus_data_30 <= __delay_data_830__delay_829_reduceadd_26 + _cond_data_23;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_834__delay_833__delay_832__delay_831__variable_11 <= __delay_data_833__delay_832__delay_831__variable_11;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_837__delay_836__delay_835_pulse_28 <= __delay_data_836__delay_835_pulse_28;
      end 
      if(_acc_1_stream_oready) begin
        _sra_data_31 <= _plus_data_30 >>> __delay_data_834__delay_833__delay_832__delay_831__variable_11;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_838__delay_837__delay_836__delay_835_pulse_28 <= __delay_data_837__delay_836__delay_835_pulse_28;
      end 
      if(__stream_conv2d_25_stream_ivalid_13 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_25 <= __delay_data_985__delay_984__delay_983____variable_281;
      end 
      if(__stream_conv2d_25_stream_ivalid_13 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_10 <= __substreamoutput_data_826;
      end 
      if(__stream_conv2d_25_stream_ivalid_13 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_11 <= __delay_data_997__delay_996__delay_995__delay_994___plus_839;
      end 
      if(__stream_conv2d_25_stream_ivalid_13 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_12 <= __delay_data_1010__delay_1009__delay_1008____variable_276;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_729 <= _acc_1_source_start;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_730 <= _tmp_729;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_731 <= _tmp_730;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_732 <= _acc_1_source_start;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_733 <= _tmp_732;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_734 <= _tmp_733;
      end 
      if(_acc_1_stream_oready && _tmp_734) begin
        __variable_wdata_25 <= 1;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_735 <= _acc_1_source_start;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_736 <= _tmp_735;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_737 <= _tmp_736;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_738 <= _tmp_737;
      end 
      if(_acc_1_stream_oready && _tmp_738) begin
        __variable_wdata_25 <= 0;
      end 
      if(_acc_1_stream_oready && 1'd0) begin
        __variable_wdata_25 <= 1;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_739 <= _acc_1_source_start;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_740 <= _tmp_739;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_741 <= _tmp_740;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_742 <= _tmp_741;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_743 <= _tmp_742;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_744 <= _tmp_743;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_745 <= _tmp_744;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_746 <= _acc_1_source_stop;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_747 <= _tmp_746;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_748 <= _tmp_747;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_749 <= _tmp_748;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_750 <= _tmp_749;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_751 <= _tmp_750;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_752 <= _tmp_751;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_753 <= _acc_1_source_busy;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_754 <= _tmp_753;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_755 <= _tmp_754;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_756 <= _tmp_755;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_757 <= _tmp_756;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_758 <= _tmp_757;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_759 <= _tmp_758;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_760 <= _acc_1_sink_busy;
      end 
      if(!_acc_1_sink_busy && _tmp_760) begin
        _acc_1_busy_reg <= 0;
      end 
      if(_acc_1_source_busy) begin
        _acc_1_busy_reg <= 1;
      end 
    end
  end

  localparam _acc_1_fsm_1 = 1;
  localparam _acc_1_fsm_2 = 2;
  localparam _acc_1_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _acc_1_fsm <= _acc_1_fsm_init;
      _acc_1_source_start <= 0;
      _acc_1_source_busy <= 0;
      _acc_1_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_25_stream_ivalid_13 && _stream_conv2d_25_stream_oready) begin
        _acc_1_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_busy) begin
        _acc_1_source_busy <= _stream_conv2d_25_source_busy;
      end 
      if(_acc_1_stream_oready && _tmp_731) begin
        _acc_1_stream_ivalid <= 1;
      end 
      if(_acc_1_stream_oready && 1'd0) begin
        _acc_1_stream_ivalid <= 0;
      end 
      case(_acc_1_fsm)
        _acc_1_fsm_init: begin
          if(_acc_1_run_flag) begin
            _acc_1_source_start <= 1;
          end 
          if(_acc_1_run_flag) begin
            _acc_1_fsm <= _acc_1_fsm_1;
          end 
        end
        _acc_1_fsm_1: begin
          if(_acc_1_source_start && _acc_1_stream_oready) begin
            _acc_1_source_start <= 0;
            _acc_1_source_busy <= 1;
          end 
          if(_acc_1_source_start && _acc_1_stream_oready) begin
            _acc_1_fsm <= _acc_1_fsm_2;
          end 
        end
        _acc_1_fsm_2: begin
          if(_acc_1_stream_oready) begin
            _acc_1_fsm <= _acc_1_fsm_3;
          end 
        end
        _acc_1_fsm_3: begin
          if(_acc_1_stream_oready && 1'd0) begin
            _acc_1_source_busy <= 0;
          end 
          if(_acc_1_stream_oready && 1'd0 && _acc_1_run_flag) begin
            _acc_1_source_start <= 1;
          end 
          if(_acc_1_stream_oready && 1'd0) begin
            _acc_1_fsm <= _acc_1_fsm_init;
          end 
          if(_acc_1_stream_oready && 1'd0 && _acc_1_run_flag) begin
            _acc_1_fsm <= _acc_1_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_2_var0_source_ram_renable <= 0;
      _add_tree_2_var0_source_fifo_deq <= 0;
      _add_tree_2_var0_idle <= 1;
      _add_tree_2_var1_source_ram_renable <= 0;
      _add_tree_2_var1_source_fifo_deq <= 0;
      _add_tree_2_var1_idle <= 1;
      _add_tree_2_var2_source_ram_renable <= 0;
      _add_tree_2_var2_source_fifo_deq <= 0;
      _add_tree_2_var2_idle <= 1;
      _add_tree_2_var3_source_ram_renable <= 0;
      _add_tree_2_var3_source_fifo_deq <= 0;
      _add_tree_2_var3_idle <= 1;
      _add_tree_2_var4_source_ram_renable <= 0;
      _add_tree_2_var4_source_fifo_deq <= 0;
      _add_tree_2_var4_idle <= 1;
      _add_tree_2_var5_source_ram_renable <= 0;
      _add_tree_2_var5_source_fifo_deq <= 0;
      _add_tree_2_var5_idle <= 1;
      _add_tree_2_var6_source_ram_renable <= 0;
      _add_tree_2_var6_source_fifo_deq <= 0;
      _add_tree_2_var6_idle <= 1;
      _add_tree_2_var7_source_ram_renable <= 0;
      _add_tree_2_var7_source_fifo_deq <= 0;
      _add_tree_2_var7_idle <= 1;
      _add_tree_2_var8_source_ram_renable <= 0;
      _add_tree_2_var8_source_fifo_deq <= 0;
      _add_tree_2_var8_idle <= 1;
      _add_tree_2_sum_sink_wenable <= 0;
      _add_tree_2_sum_sink_fifo_enq <= 0;
      __add_tree_2_stream_ivalid_1 <= 0;
      __add_tree_2_stream_ivalid_2 <= 0;
      __plusn_data_42 <= 0;
      __plusn_data_43 <= 0;
      __plusn_data_44 <= 0;
      __plusn_data_45 <= 0;
      __variable_wdata_32 <= 0;
      __variable_wdata_33 <= 0;
      __variable_wdata_34 <= 0;
      __variable_wdata_35 <= 0;
      __variable_wdata_36 <= 0;
      __variable_wdata_37 <= 0;
      __variable_wdata_38 <= 0;
      __variable_wdata_39 <= 0;
      __variable_wdata_40 <= 0;
      _tmp_713 <= 0;
      _tmp_714 <= 0;
      _tmp_715 <= 0;
      _tmp_716 <= 0;
      _tmp_717 <= 0;
      _tmp_718 <= 0;
      _tmp_719 <= 0;
      _tmp_720 <= 0;
      _tmp_721 <= 0;
      _tmp_722 <= 0;
      _tmp_723 <= 0;
      _tmp_724 <= 0;
      _tmp_725 <= 0;
      _tmp_726 <= 0;
      _tmp_727 <= 0;
      _tmp_728 <= 0;
      _add_tree_2_busy_reg <= 0;
    end else begin
      if(_add_tree_2_stream_oready) begin
        _add_tree_2_var0_source_ram_renable <= 0;
        _add_tree_2_var0_source_fifo_deq <= 0;
      end 
      _add_tree_2_var0_idle <= _add_tree_2_var0_idle;
      if(_add_tree_2_stream_oready) begin
        _add_tree_2_var1_source_ram_renable <= 0;
        _add_tree_2_var1_source_fifo_deq <= 0;
      end 
      _add_tree_2_var1_idle <= _add_tree_2_var1_idle;
      if(_add_tree_2_stream_oready) begin
        _add_tree_2_var2_source_ram_renable <= 0;
        _add_tree_2_var2_source_fifo_deq <= 0;
      end 
      _add_tree_2_var2_idle <= _add_tree_2_var2_idle;
      if(_add_tree_2_stream_oready) begin
        _add_tree_2_var3_source_ram_renable <= 0;
        _add_tree_2_var3_source_fifo_deq <= 0;
      end 
      _add_tree_2_var3_idle <= _add_tree_2_var3_idle;
      if(_add_tree_2_stream_oready) begin
        _add_tree_2_var4_source_ram_renable <= 0;
        _add_tree_2_var4_source_fifo_deq <= 0;
      end 
      _add_tree_2_var4_idle <= _add_tree_2_var4_idle;
      if(_add_tree_2_stream_oready) begin
        _add_tree_2_var5_source_ram_renable <= 0;
        _add_tree_2_var5_source_fifo_deq <= 0;
      end 
      _add_tree_2_var5_idle <= _add_tree_2_var5_idle;
      if(_add_tree_2_stream_oready) begin
        _add_tree_2_var6_source_ram_renable <= 0;
        _add_tree_2_var6_source_fifo_deq <= 0;
      end 
      _add_tree_2_var6_idle <= _add_tree_2_var6_idle;
      if(_add_tree_2_stream_oready) begin
        _add_tree_2_var7_source_ram_renable <= 0;
        _add_tree_2_var7_source_fifo_deq <= 0;
      end 
      _add_tree_2_var7_idle <= _add_tree_2_var7_idle;
      if(_add_tree_2_stream_oready) begin
        _add_tree_2_var8_source_ram_renable <= 0;
        _add_tree_2_var8_source_fifo_deq <= 0;
      end 
      _add_tree_2_var8_idle <= _add_tree_2_var8_idle;
      if(_add_tree_2_stream_oready) begin
        _add_tree_2_sum_sink_wenable <= 0;
        _add_tree_2_sum_sink_fifo_enq <= 0;
      end 
      if(_add_tree_2_stream_oready) begin
        __add_tree_2_stream_ivalid_1 <= _add_tree_2_stream_ivalid;
      end 
      if(_add_tree_2_stream_oready) begin
        __add_tree_2_stream_ivalid_2 <= __add_tree_2_stream_ivalid_1;
      end 
      if(_add_tree_2_stream_oready) begin
        __plusn_data_42 <= add_tree_2_var0_data + add_tree_2_var1_data + add_tree_2_var2_data;
      end 
      if(_add_tree_2_stream_oready) begin
        __plusn_data_43 <= add_tree_2_var3_data + add_tree_2_var4_data + add_tree_2_var5_data;
      end 
      if(_add_tree_2_stream_oready) begin
        __plusn_data_44 <= add_tree_2_var6_data + add_tree_2_var7_data + add_tree_2_var8_data;
      end 
      if(_add_tree_2_stream_oready) begin
        __plusn_data_45 <= __plusn_data_42 + __plusn_data_43 + __plusn_data_44;
      end 
      if(__stream_conv2d_25_stream_ivalid_10 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_32 <= __substreamoutput_data_672;
      end 
      if(__stream_conv2d_25_stream_ivalid_10 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_33 <= __substreamoutput_data_691;
      end 
      if(__stream_conv2d_25_stream_ivalid_10 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_34 <= __substreamoutput_data_710;
      end 
      if(__stream_conv2d_25_stream_ivalid_10 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_35 <= __substreamoutput_data_729;
      end 
      if(__stream_conv2d_25_stream_ivalid_10 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_36 <= __substreamoutput_data_748;
      end 
      if(__stream_conv2d_25_stream_ivalid_10 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_37 <= __substreamoutput_data_767;
      end 
      if(__stream_conv2d_25_stream_ivalid_10 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_38 <= __substreamoutput_data_786;
      end 
      if(__stream_conv2d_25_stream_ivalid_10 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_39 <= __substreamoutput_data_805;
      end 
      if(__stream_conv2d_25_stream_ivalid_10 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_40 <= __substreamoutput_data_824;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_713 <= _add_tree_2_source_start;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_714 <= _tmp_713;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_715 <= _tmp_714;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_716 <= _add_tree_2_source_start;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_717 <= _tmp_716;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_718 <= _tmp_717;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_719 <= _tmp_718;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_720 <= _add_tree_2_source_stop;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_721 <= _tmp_720;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_722 <= _tmp_721;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_723 <= _tmp_722;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_724 <= _add_tree_2_source_busy;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_725 <= _tmp_724;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_726 <= _tmp_725;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_727 <= _tmp_726;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_728 <= _add_tree_2_sink_busy;
      end 
      if(!_add_tree_2_sink_busy && _tmp_728) begin
        _add_tree_2_busy_reg <= 0;
      end 
      if(_add_tree_2_source_busy) begin
        _add_tree_2_busy_reg <= 1;
      end 
    end
  end

  localparam _add_tree_2_fsm_1 = 1;
  localparam _add_tree_2_fsm_2 = 2;
  localparam _add_tree_2_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_2_fsm <= _add_tree_2_fsm_init;
      _add_tree_2_source_start <= 0;
      _add_tree_2_source_busy <= 0;
      _add_tree_2_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_25_stream_ivalid_10 && _stream_conv2d_25_stream_oready) begin
        _add_tree_2_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_busy) begin
        _add_tree_2_source_busy <= _stream_conv2d_25_source_busy;
      end 
      if(_add_tree_2_stream_oready && _tmp_715) begin
        _add_tree_2_stream_ivalid <= 1;
      end 
      if(_add_tree_2_stream_oready && 1'd0) begin
        _add_tree_2_stream_ivalid <= 0;
      end 
      case(_add_tree_2_fsm)
        _add_tree_2_fsm_init: begin
          if(_add_tree_2_run_flag) begin
            _add_tree_2_source_start <= 1;
          end 
          if(_add_tree_2_run_flag) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_1;
          end 
        end
        _add_tree_2_fsm_1: begin
          if(_add_tree_2_source_start && _add_tree_2_stream_oready) begin
            _add_tree_2_source_start <= 0;
            _add_tree_2_source_busy <= 1;
          end 
          if(_add_tree_2_source_start && _add_tree_2_stream_oready) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_2;
          end 
        end
        _add_tree_2_fsm_2: begin
          if(_add_tree_2_stream_oready) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_3;
          end 
        end
        _add_tree_2_fsm_3: begin
          if(_add_tree_2_stream_oready && 1'd0) begin
            _add_tree_2_source_busy <= 0;
          end 
          if(_add_tree_2_stream_oready && 1'd0 && _add_tree_2_run_flag) begin
            _add_tree_2_source_start <= 1;
          end 
          if(_add_tree_2_stream_oready && 1'd0) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_init;
          end 
          if(_add_tree_2_stream_oready && 1'd0 && _add_tree_2_run_flag) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_round_clip_3_x_source_ram_renable <= 0;
      _mul_rshift_round_clip_3_x_source_fifo_deq <= 0;
      _mul_rshift_round_clip_3_x_idle <= 1;
      _mul_rshift_round_clip_3_y_source_ram_renable <= 0;
      _mul_rshift_round_clip_3_y_source_fifo_deq <= 0;
      _mul_rshift_round_clip_3_y_idle <= 1;
      _mul_rshift_round_clip_3_rshift_source_ram_renable <= 0;
      _mul_rshift_round_clip_3_rshift_source_fifo_deq <= 0;
      _mul_rshift_round_clip_3_rshift_idle <= 1;
      _mul_rshift_round_clip_3_z_sink_wenable <= 0;
      _mul_rshift_round_clip_3_z_sink_fifo_enq <= 0;
      __mul_rshift_round_clip_3_stream_ivalid_1 <= 0;
      __mul_rshift_round_clip_3_stream_ivalid_2 <= 0;
      __mul_rshift_round_clip_3_stream_ivalid_3 <= 0;
      __mul_rshift_round_clip_3_stream_ivalid_4 <= 0;
      __mul_rshift_round_clip_3_stream_ivalid_5 <= 0;
      __mul_rshift_round_clip_3_stream_ivalid_6 <= 0;
      __mul_rshift_round_clip_3_stream_ivalid_7 <= 0;
      __mul_rshift_round_clip_3_stream_ivalid_8 <= 0;
      _times_mul_odata_reg_49 <= 0;
      __delay_data_844_sll_55 <= 0;
      __delay_data_848__variable_48 <= 0;
      __delay_data_852_eq_67 <= 0;
      __delay_data_845__delay_844_sll_55 <= 0;
      __delay_data_849__delay_848__variable_48 <= 0;
      __delay_data_853__delay_852_eq_67 <= 0;
      __delay_data_846__delay_845__delay_844_sll_55 <= 0;
      __delay_data_850__delay_849__delay_848__variable_48 <= 0;
      __delay_data_854__delay_853__delay_852_eq_67 <= 0;
      __delay_data_847__delay_846__delay_845__delay_844_sll_55 <= 0;
      __delay_data_851__delay_850__delay_849__delay_848__variable_48 <= 0;
      __delay_data_855__delay_854__delay_853__delay_852_eq_67 <= 0;
      _cond_data_68 <= 0;
      _greaterthan_data_69 <= 0;
      _lessthan_data_73 <= 0;
      _greatereq_data_77 <= 0;
      __delay_data_856_cond_68 <= 0;
      _cond_data_71 <= 0;
      _cond_data_75 <= 0;
      __delay_data_857_greatereq_77 <= 0;
      _cond_data_79 <= 0;
      __variable_wdata_46 <= 0;
      __variable_wdata_47 <= 0;
      __variable_wdata_48 <= 0;
      _tmp_761 <= 0;
      _tmp_762 <= 0;
      _tmp_763 <= 0;
      _tmp_764 <= 0;
      _tmp_765 <= 0;
      _tmp_766 <= 0;
      _tmp_767 <= 0;
      _tmp_768 <= 0;
      _tmp_769 <= 0;
      _tmp_770 <= 0;
      _tmp_771 <= 0;
      _tmp_772 <= 0;
      _tmp_773 <= 0;
      _tmp_774 <= 0;
      _tmp_775 <= 0;
      _tmp_776 <= 0;
      _tmp_777 <= 0;
      _tmp_778 <= 0;
      _tmp_779 <= 0;
      _tmp_780 <= 0;
      _tmp_781 <= 0;
      _tmp_782 <= 0;
      _tmp_783 <= 0;
      _tmp_784 <= 0;
      _tmp_785 <= 0;
      _tmp_786 <= 0;
      _tmp_787 <= 0;
      _tmp_788 <= 0;
      _tmp_789 <= 0;
      _tmp_790 <= 0;
      _tmp_791 <= 0;
      _tmp_792 <= 0;
      _tmp_793 <= 0;
      _tmp_794 <= 0;
      _mul_rshift_round_clip_3_busy_reg <= 0;
    end else begin
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _mul_rshift_round_clip_3_x_source_ram_renable <= 0;
        _mul_rshift_round_clip_3_x_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_3_x_idle <= _mul_rshift_round_clip_3_x_idle;
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _mul_rshift_round_clip_3_y_source_ram_renable <= 0;
        _mul_rshift_round_clip_3_y_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_3_y_idle <= _mul_rshift_round_clip_3_y_idle;
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _mul_rshift_round_clip_3_rshift_source_ram_renable <= 0;
        _mul_rshift_round_clip_3_rshift_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_3_rshift_idle <= _mul_rshift_round_clip_3_rshift_idle;
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _mul_rshift_round_clip_3_z_sink_wenable <= 0;
        _mul_rshift_round_clip_3_z_sink_fifo_enq <= 0;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __mul_rshift_round_clip_3_stream_ivalid_1 <= _mul_rshift_round_clip_3_stream_ivalid;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __mul_rshift_round_clip_3_stream_ivalid_2 <= __mul_rshift_round_clip_3_stream_ivalid_1;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __mul_rshift_round_clip_3_stream_ivalid_3 <= __mul_rshift_round_clip_3_stream_ivalid_2;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __mul_rshift_round_clip_3_stream_ivalid_4 <= __mul_rshift_round_clip_3_stream_ivalid_3;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __mul_rshift_round_clip_3_stream_ivalid_5 <= __mul_rshift_round_clip_3_stream_ivalid_4;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __mul_rshift_round_clip_3_stream_ivalid_6 <= __mul_rshift_round_clip_3_stream_ivalid_5;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __mul_rshift_round_clip_3_stream_ivalid_7 <= __mul_rshift_round_clip_3_stream_ivalid_6;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __mul_rshift_round_clip_3_stream_ivalid_8 <= __mul_rshift_round_clip_3_stream_ivalid_7;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _times_mul_odata_reg_49 <= _times_mul_odata_49;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __delay_data_844_sll_55 <= _sll_data_55;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __delay_data_848__variable_48 <= mul_rshift_round_clip_3_rshift_data;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __delay_data_852_eq_67 <= _eq_data_67;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __delay_data_845__delay_844_sll_55 <= __delay_data_844_sll_55;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __delay_data_849__delay_848__variable_48 <= __delay_data_848__variable_48;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __delay_data_853__delay_852_eq_67 <= __delay_data_852_eq_67;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __delay_data_846__delay_845__delay_844_sll_55 <= __delay_data_845__delay_844_sll_55;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __delay_data_850__delay_849__delay_848__variable_48 <= __delay_data_849__delay_848__variable_48;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __delay_data_854__delay_853__delay_852_eq_67 <= __delay_data_853__delay_852_eq_67;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __delay_data_847__delay_846__delay_845__delay_844_sll_55 <= __delay_data_846__delay_845__delay_844_sll_55;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __delay_data_851__delay_850__delay_849__delay_848__variable_48 <= __delay_data_850__delay_849__delay_848__variable_48;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __delay_data_855__delay_854__delay_853__delay_852_eq_67 <= __delay_data_854__delay_853__delay_852_eq_67;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _cond_data_68 <= (__delay_data_855__delay_854__delay_853__delay_852_eq_67)? _times_data_49 : _sra_data_65;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _greaterthan_data_69 <= _cond_data_68 > 32'sd2147483647;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _lessthan_data_73 <= _cond_data_68 < -32'sd2147483647;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _greatereq_data_77 <= _cond_data_68 >= 1'sd0;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __delay_data_856_cond_68 <= _cond_data_68;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _cond_data_71 <= (_greaterthan_data_69)? 32'sd2147483647 : __delay_data_856_cond_68;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _cond_data_75 <= (_lessthan_data_73)? -32'sd2147483647 : __delay_data_856_cond_68;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        __delay_data_857_greatereq_77 <= _greatereq_data_77;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _cond_data_79 <= (__delay_data_857_greatereq_77)? _cond_data_71 : _cond_data_75;
      end 
      if(__stream_conv2d_25_stream_ivalid_20 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_46 <= _plus_data_842;
      end 
      if(__stream_conv2d_25_stream_ivalid_20 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_47 <= __delay_data_1049__delay_1048__delay_1047__delay_1046___cond_304;
      end 
      if(__stream_conv2d_25_stream_ivalid_20 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_48 <= __delay_data_1068__delay_1067__delay_1066__delay_1065___plus_858;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_761 <= _mul_rshift_round_clip_3_source_start;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_762 <= _tmp_761;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_763 <= _tmp_762;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_764 <= _mul_rshift_round_clip_3_source_start;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_765 <= _tmp_764;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_766 <= _tmp_765;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_767 <= _tmp_766;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_768 <= _tmp_767;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_769 <= _tmp_768;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_770 <= _tmp_769;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_771 <= _tmp_770;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_772 <= _tmp_771;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_773 <= _tmp_772;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_774 <= _mul_rshift_round_clip_3_source_stop;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_775 <= _tmp_774;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_776 <= _tmp_775;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_777 <= _tmp_776;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_778 <= _tmp_777;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_779 <= _tmp_778;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_780 <= _tmp_779;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_781 <= _tmp_780;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_782 <= _tmp_781;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_783 <= _tmp_782;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_784 <= _mul_rshift_round_clip_3_source_busy;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_785 <= _tmp_784;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_786 <= _tmp_785;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_787 <= _tmp_786;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_788 <= _tmp_787;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_789 <= _tmp_788;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_790 <= _tmp_789;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_791 <= _tmp_790;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_792 <= _tmp_791;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_793 <= _tmp_792;
      end 
      if(_mul_rshift_round_clip_3_stream_oready) begin
        _tmp_794 <= _mul_rshift_round_clip_3_sink_busy;
      end 
      if(!_mul_rshift_round_clip_3_sink_busy && _tmp_794) begin
        _mul_rshift_round_clip_3_busy_reg <= 0;
      end 
      if(_mul_rshift_round_clip_3_source_busy) begin
        _mul_rshift_round_clip_3_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_rshift_round_clip_3_fsm_1 = 1;
  localparam _mul_rshift_round_clip_3_fsm_2 = 2;
  localparam _mul_rshift_round_clip_3_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_round_clip_3_fsm <= _mul_rshift_round_clip_3_fsm_init;
      _mul_rshift_round_clip_3_source_start <= 0;
      _mul_rshift_round_clip_3_source_busy <= 0;
      _mul_rshift_round_clip_3_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_25_stream_ivalid_20 && _stream_conv2d_25_stream_oready) begin
        _mul_rshift_round_clip_3_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_busy) begin
        _mul_rshift_round_clip_3_source_busy <= _stream_conv2d_25_source_busy;
      end 
      if(_mul_rshift_round_clip_3_stream_oready && _tmp_763) begin
        _mul_rshift_round_clip_3_stream_ivalid <= 1;
      end 
      if(_mul_rshift_round_clip_3_stream_oready && 1'd0) begin
        _mul_rshift_round_clip_3_stream_ivalid <= 0;
      end 
      case(_mul_rshift_round_clip_3_fsm)
        _mul_rshift_round_clip_3_fsm_init: begin
          if(_mul_rshift_round_clip_3_run_flag) begin
            _mul_rshift_round_clip_3_source_start <= 1;
          end 
          if(_mul_rshift_round_clip_3_run_flag) begin
            _mul_rshift_round_clip_3_fsm <= _mul_rshift_round_clip_3_fsm_1;
          end 
        end
        _mul_rshift_round_clip_3_fsm_1: begin
          if(_mul_rshift_round_clip_3_source_start && _mul_rshift_round_clip_3_stream_oready) begin
            _mul_rshift_round_clip_3_source_start <= 0;
            _mul_rshift_round_clip_3_source_busy <= 1;
          end 
          if(_mul_rshift_round_clip_3_source_start && _mul_rshift_round_clip_3_stream_oready) begin
            _mul_rshift_round_clip_3_fsm <= _mul_rshift_round_clip_3_fsm_2;
          end 
        end
        _mul_rshift_round_clip_3_fsm_2: begin
          if(_mul_rshift_round_clip_3_stream_oready) begin
            _mul_rshift_round_clip_3_fsm <= _mul_rshift_round_clip_3_fsm_3;
          end 
        end
        _mul_rshift_round_clip_3_fsm_3: begin
          if(_mul_rshift_round_clip_3_stream_oready && 1'd0) begin
            _mul_rshift_round_clip_3_source_busy <= 0;
          end 
          if(_mul_rshift_round_clip_3_stream_oready && 1'd0 && _mul_rshift_round_clip_3_run_flag) begin
            _mul_rshift_round_clip_3_source_start <= 1;
          end 
          if(_mul_rshift_round_clip_3_stream_oready && 1'd0) begin
            _mul_rshift_round_clip_3_fsm <= _mul_rshift_round_clip_3_fsm_init;
          end 
          if(_mul_rshift_round_clip_3_stream_oready && 1'd0 && _mul_rshift_round_clip_3_run_flag) begin
            _mul_rshift_round_clip_3_fsm <= _mul_rshift_round_clip_3_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_4_x_source_ram_renable <= 0;
      _mul_4_x_source_fifo_deq <= 0;
      _mul_4_x_idle <= 1;
      _mul_4_y_source_ram_renable <= 0;
      _mul_4_y_source_fifo_deq <= 0;
      _mul_4_y_idle <= 1;
      _mul_4_rshift_source_ram_renable <= 0;
      _mul_4_rshift_source_fifo_deq <= 0;
      _mul_4_rshift_idle <= 1;
      _mul_4_z_sink_wenable <= 0;
      _mul_4_z_sink_fifo_enq <= 0;
      __mul_4_stream_ivalid_1 <= 0;
      __mul_4_stream_ivalid_2 <= 0;
      __mul_4_stream_ivalid_3 <= 0;
      __mul_4_stream_ivalid_4 <= 0;
      __mul_4_stream_ivalid_5 <= 0;
      __mul_4_stream_ivalid_6 <= 0;
      __mul_4_stream_ivalid_7 <= 0;
      __mul_4_stream_ivalid_8 <= 0;
      _greaterthan_data_83 <= 0;
      _minus_data_85 <= 0;
      _greatereq_data_96 <= 0;
      __delay_data_658__variable_80 <= 0;
      __delay_data_661__variable_81 <= 0;
      __delay_data_664__variable_82 <= 0;
      _sll_data_87 <= 0;
      __delay_data_655_greaterthan_83 <= 0;
      __delay_data_656_greatereq_96 <= 0;
      __delay_data_659__delay_658__variable_80 <= 0;
      __delay_data_662__delay_661__variable_81 <= 0;
      __delay_data_665__delay_664__variable_82 <= 0;
      _cond_data_93 <= 0;
      __delay_data_657__delay_656_greatereq_96 <= 0;
      __delay_data_660__delay_659__delay_658__variable_80 <= 0;
      __delay_data_663__delay_662__delay_661__variable_81 <= 0;
      __delay_data_666__delay_665__delay_664__variable_82 <= 0;
      __muladd_madd_odata_reg_99 <= 0;
      __delay_data_667__delay_666__delay_665__delay_664__variable_82 <= 0;
      __delay_data_668__delay_667__delay_666__delay_665____variable_82 <= 0;
      __delay_data_669__delay_668__delay_667__delay_666____variable_82 <= 0;
      __delay_data_670__delay_669__delay_668__delay_667____variable_82 <= 0;
      _sra_data_100 <= 0;
      __variable_wdata_80 <= 0;
      __variable_wdata_81 <= 0;
      __variable_wdata_82 <= 0;
      _tmp_407 <= 0;
      _tmp_408 <= 0;
      _tmp_409 <= 0;
      _tmp_410 <= 0;
      _tmp_411 <= 0;
      _tmp_412 <= 0;
      _tmp_413 <= 0;
      _tmp_414 <= 0;
      _tmp_415 <= 0;
      _tmp_416 <= 0;
      _tmp_417 <= 0;
      _tmp_418 <= 0;
      _tmp_419 <= 0;
      _tmp_420 <= 0;
      _tmp_421 <= 0;
      _tmp_422 <= 0;
      _tmp_423 <= 0;
      _tmp_424 <= 0;
      _tmp_425 <= 0;
      _tmp_426 <= 0;
      _tmp_427 <= 0;
      _tmp_428 <= 0;
      _tmp_429 <= 0;
      _tmp_430 <= 0;
      _tmp_431 <= 0;
      _tmp_432 <= 0;
      _tmp_433 <= 0;
      _tmp_434 <= 0;
      _tmp_435 <= 0;
      _tmp_436 <= 0;
      _tmp_437 <= 0;
      _tmp_438 <= 0;
      _tmp_439 <= 0;
      _tmp_440 <= 0;
      _mul_4_busy_reg <= 0;
    end else begin
      if(_mul_4_stream_oready) begin
        _mul_4_x_source_ram_renable <= 0;
        _mul_4_x_source_fifo_deq <= 0;
      end 
      _mul_4_x_idle <= _mul_4_x_idle;
      if(_mul_4_stream_oready) begin
        _mul_4_y_source_ram_renable <= 0;
        _mul_4_y_source_fifo_deq <= 0;
      end 
      _mul_4_y_idle <= _mul_4_y_idle;
      if(_mul_4_stream_oready) begin
        _mul_4_rshift_source_ram_renable <= 0;
        _mul_4_rshift_source_fifo_deq <= 0;
      end 
      _mul_4_rshift_idle <= _mul_4_rshift_idle;
      if(_mul_4_stream_oready) begin
        _mul_4_z_sink_wenable <= 0;
        _mul_4_z_sink_fifo_enq <= 0;
      end 
      if(_mul_4_stream_oready) begin
        __mul_4_stream_ivalid_1 <= _mul_4_stream_ivalid;
      end 
      if(_mul_4_stream_oready) begin
        __mul_4_stream_ivalid_2 <= __mul_4_stream_ivalid_1;
      end 
      if(_mul_4_stream_oready) begin
        __mul_4_stream_ivalid_3 <= __mul_4_stream_ivalid_2;
      end 
      if(_mul_4_stream_oready) begin
        __mul_4_stream_ivalid_4 <= __mul_4_stream_ivalid_3;
      end 
      if(_mul_4_stream_oready) begin
        __mul_4_stream_ivalid_5 <= __mul_4_stream_ivalid_4;
      end 
      if(_mul_4_stream_oready) begin
        __mul_4_stream_ivalid_6 <= __mul_4_stream_ivalid_5;
      end 
      if(_mul_4_stream_oready) begin
        __mul_4_stream_ivalid_7 <= __mul_4_stream_ivalid_6;
      end 
      if(_mul_4_stream_oready) begin
        __mul_4_stream_ivalid_8 <= __mul_4_stream_ivalid_7;
      end 
      if(_mul_4_stream_oready) begin
        _greaterthan_data_83 <= mul_4_rshift_data > 1'sd0;
      end 
      if(_mul_4_stream_oready) begin
        _minus_data_85 <= mul_4_rshift_data - 2'sd1;
      end 
      if(_mul_4_stream_oready) begin
        _greatereq_data_96 <= mul_4_x_data >= 1'sd0;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_658__variable_80 <= mul_4_x_data;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_661__variable_81 <= mul_4_y_data;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_664__variable_82 <= mul_4_rshift_data;
      end 
      if(_mul_4_stream_oready) begin
        _sll_data_87 <= 2'sd1 << _minus_data_85;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_655_greaterthan_83 <= _greaterthan_data_83;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_656_greatereq_96 <= _greatereq_data_96;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_659__delay_658__variable_80 <= __delay_data_658__variable_80;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_662__delay_661__variable_81 <= __delay_data_661__variable_81;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_665__delay_664__variable_82 <= __delay_data_664__variable_82;
      end 
      if(_mul_4_stream_oready) begin
        _cond_data_93 <= (__delay_data_655_greaterthan_83)? _sll_data_87 : 1'sd0;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_657__delay_656_greatereq_96 <= __delay_data_656_greatereq_96;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_660__delay_659__delay_658__variable_80 <= __delay_data_659__delay_658__variable_80;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_663__delay_662__delay_661__variable_81 <= __delay_data_662__delay_661__variable_81;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_666__delay_665__delay_664__variable_82 <= __delay_data_665__delay_664__variable_82;
      end 
      if(_mul_4_stream_oready) begin
        __muladd_madd_odata_reg_99 <= __muladd_madd_odata_99;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_667__delay_666__delay_665__delay_664__variable_82 <= __delay_data_666__delay_665__delay_664__variable_82;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_668__delay_667__delay_666__delay_665____variable_82 <= __delay_data_667__delay_666__delay_665__delay_664__variable_82;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_669__delay_668__delay_667__delay_666____variable_82 <= __delay_data_668__delay_667__delay_666__delay_665____variable_82;
      end 
      if(_mul_4_stream_oready) begin
        __delay_data_670__delay_669__delay_668__delay_667____variable_82 <= __delay_data_669__delay_668__delay_667__delay_666____variable_82;
      end 
      if(_mul_4_stream_oready) begin
        _sra_data_100 <= __muladd_data_99 >>> __delay_data_670__delay_669__delay_668__delay_667____variable_82;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_80 <= _cond_data_637;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_81 <= __delay_data_956_reinterpretcast_609;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_82 <= _plus_data_671;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_407 <= _mul_4_source_start;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_408 <= _tmp_407;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_409 <= _tmp_408;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_410 <= _mul_4_source_start;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_411 <= _tmp_410;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_412 <= _tmp_411;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_413 <= _tmp_412;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_414 <= _tmp_413;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_415 <= _tmp_414;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_416 <= _tmp_415;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_417 <= _tmp_416;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_418 <= _tmp_417;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_419 <= _tmp_418;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_420 <= _mul_4_source_stop;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_421 <= _tmp_420;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_422 <= _tmp_421;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_423 <= _tmp_422;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_424 <= _tmp_423;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_425 <= _tmp_424;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_426 <= _tmp_425;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_427 <= _tmp_426;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_428 <= _tmp_427;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_429 <= _tmp_428;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_430 <= _mul_4_source_busy;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_431 <= _tmp_430;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_432 <= _tmp_431;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_433 <= _tmp_432;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_434 <= _tmp_433;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_435 <= _tmp_434;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_436 <= _tmp_435;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_437 <= _tmp_436;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_438 <= _tmp_437;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_439 <= _tmp_438;
      end 
      if(_mul_4_stream_oready) begin
        _tmp_440 <= _mul_4_sink_busy;
      end 
      if(!_mul_4_sink_busy && _tmp_440) begin
        _mul_4_busy_reg <= 0;
      end 
      if(_mul_4_source_busy) begin
        _mul_4_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_4_fsm_1 = 1;
  localparam _mul_4_fsm_2 = 2;
  localparam _mul_4_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_4_fsm <= _mul_4_fsm_init;
      _mul_4_source_start <= 0;
      _mul_4_source_busy <= 0;
      _mul_4_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        _mul_4_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_busy) begin
        _mul_4_source_busy <= _stream_conv2d_25_source_busy;
      end 
      if(_mul_4_stream_oready && _tmp_409) begin
        _mul_4_stream_ivalid <= 1;
      end 
      if(_mul_4_stream_oready && 1'd0) begin
        _mul_4_stream_ivalid <= 0;
      end 
      case(_mul_4_fsm)
        _mul_4_fsm_init: begin
          if(_mul_4_run_flag) begin
            _mul_4_source_start <= 1;
          end 
          if(_mul_4_run_flag) begin
            _mul_4_fsm <= _mul_4_fsm_1;
          end 
        end
        _mul_4_fsm_1: begin
          if(_mul_4_source_start && _mul_4_stream_oready) begin
            _mul_4_source_start <= 0;
            _mul_4_source_busy <= 1;
          end 
          if(_mul_4_source_start && _mul_4_stream_oready) begin
            _mul_4_fsm <= _mul_4_fsm_2;
          end 
        end
        _mul_4_fsm_2: begin
          if(_mul_4_stream_oready) begin
            _mul_4_fsm <= _mul_4_fsm_3;
          end 
        end
        _mul_4_fsm_3: begin
          if(_mul_4_stream_oready && 1'd0) begin
            _mul_4_source_busy <= 0;
          end 
          if(_mul_4_stream_oready && 1'd0 && _mul_4_run_flag) begin
            _mul_4_source_start <= 1;
          end 
          if(_mul_4_stream_oready && 1'd0) begin
            _mul_4_fsm <= _mul_4_fsm_init;
          end 
          if(_mul_4_stream_oready && 1'd0 && _mul_4_run_flag) begin
            _mul_4_fsm <= _mul_4_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_5_x_source_ram_renable <= 0;
      _mul_5_x_source_fifo_deq <= 0;
      _mul_5_x_idle <= 1;
      _mul_5_y_source_ram_renable <= 0;
      _mul_5_y_source_fifo_deq <= 0;
      _mul_5_y_idle <= 1;
      _mul_5_rshift_source_ram_renable <= 0;
      _mul_5_rshift_source_fifo_deq <= 0;
      _mul_5_rshift_idle <= 1;
      _mul_5_z_sink_wenable <= 0;
      _mul_5_z_sink_fifo_enq <= 0;
      __mul_5_stream_ivalid_1 <= 0;
      __mul_5_stream_ivalid_2 <= 0;
      __mul_5_stream_ivalid_3 <= 0;
      __mul_5_stream_ivalid_4 <= 0;
      __mul_5_stream_ivalid_5 <= 0;
      __mul_5_stream_ivalid_6 <= 0;
      __mul_5_stream_ivalid_7 <= 0;
      __mul_5_stream_ivalid_8 <= 0;
      _greaterthan_data_104 <= 0;
      _minus_data_106 <= 0;
      _greatereq_data_117 <= 0;
      __delay_data_677__variable_101 <= 0;
      __delay_data_680__variable_102 <= 0;
      __delay_data_683__variable_103 <= 0;
      _sll_data_108 <= 0;
      __delay_data_674_greaterthan_104 <= 0;
      __delay_data_675_greatereq_117 <= 0;
      __delay_data_678__delay_677__variable_101 <= 0;
      __delay_data_681__delay_680__variable_102 <= 0;
      __delay_data_684__delay_683__variable_103 <= 0;
      _cond_data_114 <= 0;
      __delay_data_676__delay_675_greatereq_117 <= 0;
      __delay_data_679__delay_678__delay_677__variable_101 <= 0;
      __delay_data_682__delay_681__delay_680__variable_102 <= 0;
      __delay_data_685__delay_684__delay_683__variable_103 <= 0;
      __muladd_madd_odata_reg_120 <= 0;
      __delay_data_686__delay_685__delay_684____variable_103 <= 0;
      __delay_data_687__delay_686__delay_685____variable_103 <= 0;
      __delay_data_688__delay_687__delay_686____variable_103 <= 0;
      __delay_data_689__delay_688__delay_687____variable_103 <= 0;
      _sra_data_121 <= 0;
      __variable_wdata_101 <= 0;
      __variable_wdata_102 <= 0;
      __variable_wdata_103 <= 0;
      _tmp_441 <= 0;
      _tmp_442 <= 0;
      _tmp_443 <= 0;
      _tmp_444 <= 0;
      _tmp_445 <= 0;
      _tmp_446 <= 0;
      _tmp_447 <= 0;
      _tmp_448 <= 0;
      _tmp_449 <= 0;
      _tmp_450 <= 0;
      _tmp_451 <= 0;
      _tmp_452 <= 0;
      _tmp_453 <= 0;
      _tmp_454 <= 0;
      _tmp_455 <= 0;
      _tmp_456 <= 0;
      _tmp_457 <= 0;
      _tmp_458 <= 0;
      _tmp_459 <= 0;
      _tmp_460 <= 0;
      _tmp_461 <= 0;
      _tmp_462 <= 0;
      _tmp_463 <= 0;
      _tmp_464 <= 0;
      _tmp_465 <= 0;
      _tmp_466 <= 0;
      _tmp_467 <= 0;
      _tmp_468 <= 0;
      _tmp_469 <= 0;
      _tmp_470 <= 0;
      _tmp_471 <= 0;
      _tmp_472 <= 0;
      _tmp_473 <= 0;
      _tmp_474 <= 0;
      _mul_5_busy_reg <= 0;
    end else begin
      if(_mul_5_stream_oready) begin
        _mul_5_x_source_ram_renable <= 0;
        _mul_5_x_source_fifo_deq <= 0;
      end 
      _mul_5_x_idle <= _mul_5_x_idle;
      if(_mul_5_stream_oready) begin
        _mul_5_y_source_ram_renable <= 0;
        _mul_5_y_source_fifo_deq <= 0;
      end 
      _mul_5_y_idle <= _mul_5_y_idle;
      if(_mul_5_stream_oready) begin
        _mul_5_rshift_source_ram_renable <= 0;
        _mul_5_rshift_source_fifo_deq <= 0;
      end 
      _mul_5_rshift_idle <= _mul_5_rshift_idle;
      if(_mul_5_stream_oready) begin
        _mul_5_z_sink_wenable <= 0;
        _mul_5_z_sink_fifo_enq <= 0;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_1 <= _mul_5_stream_ivalid;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_2 <= __mul_5_stream_ivalid_1;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_3 <= __mul_5_stream_ivalid_2;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_4 <= __mul_5_stream_ivalid_3;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_5 <= __mul_5_stream_ivalid_4;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_6 <= __mul_5_stream_ivalid_5;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_7 <= __mul_5_stream_ivalid_6;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_8 <= __mul_5_stream_ivalid_7;
      end 
      if(_mul_5_stream_oready) begin
        _greaterthan_data_104 <= mul_5_rshift_data > 1'sd0;
      end 
      if(_mul_5_stream_oready) begin
        _minus_data_106 <= mul_5_rshift_data - 2'sd1;
      end 
      if(_mul_5_stream_oready) begin
        _greatereq_data_117 <= mul_5_x_data >= 1'sd0;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_677__variable_101 <= mul_5_x_data;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_680__variable_102 <= mul_5_y_data;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_683__variable_103 <= mul_5_rshift_data;
      end 
      if(_mul_5_stream_oready) begin
        _sll_data_108 <= 2'sd1 << _minus_data_106;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_674_greaterthan_104 <= _greaterthan_data_104;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_675_greatereq_117 <= _greatereq_data_117;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_678__delay_677__variable_101 <= __delay_data_677__variable_101;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_681__delay_680__variable_102 <= __delay_data_680__variable_102;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_684__delay_683__variable_103 <= __delay_data_683__variable_103;
      end 
      if(_mul_5_stream_oready) begin
        _cond_data_114 <= (__delay_data_674_greaterthan_104)? _sll_data_108 : 1'sd0;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_676__delay_675_greatereq_117 <= __delay_data_675_greatereq_117;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_679__delay_678__delay_677__variable_101 <= __delay_data_678__delay_677__variable_101;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_682__delay_681__delay_680__variable_102 <= __delay_data_681__delay_680__variable_102;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_685__delay_684__delay_683__variable_103 <= __delay_data_684__delay_683__variable_103;
      end 
      if(_mul_5_stream_oready) begin
        __muladd_madd_odata_reg_120 <= __muladd_madd_odata_120;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_686__delay_685__delay_684____variable_103 <= __delay_data_685__delay_684__delay_683__variable_103;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_687__delay_686__delay_685____variable_103 <= __delay_data_686__delay_685__delay_684____variable_103;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_688__delay_687__delay_686____variable_103 <= __delay_data_687__delay_686__delay_685____variable_103;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_689__delay_688__delay_687____variable_103 <= __delay_data_688__delay_687__delay_686____variable_103;
      end 
      if(_mul_5_stream_oready) begin
        _sra_data_121 <= __muladd_data_120 >>> __delay_data_689__delay_688__delay_687____variable_103;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_101 <= _cond_data_639;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_102 <= __delay_data_958_reinterpretcast_610;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_103 <= _plus_data_690;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_441 <= _mul_5_source_start;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_442 <= _tmp_441;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_443 <= _tmp_442;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_444 <= _mul_5_source_start;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_445 <= _tmp_444;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_446 <= _tmp_445;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_447 <= _tmp_446;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_448 <= _tmp_447;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_449 <= _tmp_448;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_450 <= _tmp_449;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_451 <= _tmp_450;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_452 <= _tmp_451;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_453 <= _tmp_452;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_454 <= _mul_5_source_stop;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_455 <= _tmp_454;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_456 <= _tmp_455;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_457 <= _tmp_456;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_458 <= _tmp_457;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_459 <= _tmp_458;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_460 <= _tmp_459;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_461 <= _tmp_460;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_462 <= _tmp_461;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_463 <= _tmp_462;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_464 <= _mul_5_source_busy;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_465 <= _tmp_464;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_466 <= _tmp_465;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_467 <= _tmp_466;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_468 <= _tmp_467;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_469 <= _tmp_468;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_470 <= _tmp_469;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_471 <= _tmp_470;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_472 <= _tmp_471;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_473 <= _tmp_472;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_474 <= _mul_5_sink_busy;
      end 
      if(!_mul_5_sink_busy && _tmp_474) begin
        _mul_5_busy_reg <= 0;
      end 
      if(_mul_5_source_busy) begin
        _mul_5_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_5_fsm_1 = 1;
  localparam _mul_5_fsm_2 = 2;
  localparam _mul_5_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_5_fsm <= _mul_5_fsm_init;
      _mul_5_source_start <= 0;
      _mul_5_source_busy <= 0;
      _mul_5_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        _mul_5_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_busy) begin
        _mul_5_source_busy <= _stream_conv2d_25_source_busy;
      end 
      if(_mul_5_stream_oready && _tmp_443) begin
        _mul_5_stream_ivalid <= 1;
      end 
      if(_mul_5_stream_oready && 1'd0) begin
        _mul_5_stream_ivalid <= 0;
      end 
      case(_mul_5_fsm)
        _mul_5_fsm_init: begin
          if(_mul_5_run_flag) begin
            _mul_5_source_start <= 1;
          end 
          if(_mul_5_run_flag) begin
            _mul_5_fsm <= _mul_5_fsm_1;
          end 
        end
        _mul_5_fsm_1: begin
          if(_mul_5_source_start && _mul_5_stream_oready) begin
            _mul_5_source_start <= 0;
            _mul_5_source_busy <= 1;
          end 
          if(_mul_5_source_start && _mul_5_stream_oready) begin
            _mul_5_fsm <= _mul_5_fsm_2;
          end 
        end
        _mul_5_fsm_2: begin
          if(_mul_5_stream_oready) begin
            _mul_5_fsm <= _mul_5_fsm_3;
          end 
        end
        _mul_5_fsm_3: begin
          if(_mul_5_stream_oready && 1'd0) begin
            _mul_5_source_busy <= 0;
          end 
          if(_mul_5_stream_oready && 1'd0 && _mul_5_run_flag) begin
            _mul_5_source_start <= 1;
          end 
          if(_mul_5_stream_oready && 1'd0) begin
            _mul_5_fsm <= _mul_5_fsm_init;
          end 
          if(_mul_5_stream_oready && 1'd0 && _mul_5_run_flag) begin
            _mul_5_fsm <= _mul_5_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_6_x_source_ram_renable <= 0;
      _mul_6_x_source_fifo_deq <= 0;
      _mul_6_x_idle <= 1;
      _mul_6_y_source_ram_renable <= 0;
      _mul_6_y_source_fifo_deq <= 0;
      _mul_6_y_idle <= 1;
      _mul_6_rshift_source_ram_renable <= 0;
      _mul_6_rshift_source_fifo_deq <= 0;
      _mul_6_rshift_idle <= 1;
      _mul_6_z_sink_wenable <= 0;
      _mul_6_z_sink_fifo_enq <= 0;
      __mul_6_stream_ivalid_1 <= 0;
      __mul_6_stream_ivalid_2 <= 0;
      __mul_6_stream_ivalid_3 <= 0;
      __mul_6_stream_ivalid_4 <= 0;
      __mul_6_stream_ivalid_5 <= 0;
      __mul_6_stream_ivalid_6 <= 0;
      __mul_6_stream_ivalid_7 <= 0;
      __mul_6_stream_ivalid_8 <= 0;
      _greaterthan_data_125 <= 0;
      _minus_data_127 <= 0;
      _greatereq_data_138 <= 0;
      __delay_data_696__variable_122 <= 0;
      __delay_data_699__variable_123 <= 0;
      __delay_data_702__variable_124 <= 0;
      _sll_data_129 <= 0;
      __delay_data_693_greaterthan_125 <= 0;
      __delay_data_694_greatereq_138 <= 0;
      __delay_data_697__delay_696__variable_122 <= 0;
      __delay_data_700__delay_699__variable_123 <= 0;
      __delay_data_703__delay_702__variable_124 <= 0;
      _cond_data_135 <= 0;
      __delay_data_695__delay_694_greatereq_138 <= 0;
      __delay_data_698__delay_697__delay_696__variable_122 <= 0;
      __delay_data_701__delay_700__delay_699__variable_123 <= 0;
      __delay_data_704__delay_703__delay_702__variable_124 <= 0;
      __muladd_madd_odata_reg_141 <= 0;
      __delay_data_705__delay_704__delay_703____variable_124 <= 0;
      __delay_data_706__delay_705__delay_704____variable_124 <= 0;
      __delay_data_707__delay_706__delay_705____variable_124 <= 0;
      __delay_data_708__delay_707__delay_706____variable_124 <= 0;
      _sra_data_142 <= 0;
      __variable_wdata_122 <= 0;
      __variable_wdata_123 <= 0;
      __variable_wdata_124 <= 0;
      _tmp_475 <= 0;
      _tmp_476 <= 0;
      _tmp_477 <= 0;
      _tmp_478 <= 0;
      _tmp_479 <= 0;
      _tmp_480 <= 0;
      _tmp_481 <= 0;
      _tmp_482 <= 0;
      _tmp_483 <= 0;
      _tmp_484 <= 0;
      _tmp_485 <= 0;
      _tmp_486 <= 0;
      _tmp_487 <= 0;
      _tmp_488 <= 0;
      _tmp_489 <= 0;
      _tmp_490 <= 0;
      _tmp_491 <= 0;
      _tmp_492 <= 0;
      _tmp_493 <= 0;
      _tmp_494 <= 0;
      _tmp_495 <= 0;
      _tmp_496 <= 0;
      _tmp_497 <= 0;
      _tmp_498 <= 0;
      _tmp_499 <= 0;
      _tmp_500 <= 0;
      _tmp_501 <= 0;
      _tmp_502 <= 0;
      _tmp_503 <= 0;
      _tmp_504 <= 0;
      _tmp_505 <= 0;
      _tmp_506 <= 0;
      _tmp_507 <= 0;
      _tmp_508 <= 0;
      _mul_6_busy_reg <= 0;
    end else begin
      if(_mul_6_stream_oready) begin
        _mul_6_x_source_ram_renable <= 0;
        _mul_6_x_source_fifo_deq <= 0;
      end 
      _mul_6_x_idle <= _mul_6_x_idle;
      if(_mul_6_stream_oready) begin
        _mul_6_y_source_ram_renable <= 0;
        _mul_6_y_source_fifo_deq <= 0;
      end 
      _mul_6_y_idle <= _mul_6_y_idle;
      if(_mul_6_stream_oready) begin
        _mul_6_rshift_source_ram_renable <= 0;
        _mul_6_rshift_source_fifo_deq <= 0;
      end 
      _mul_6_rshift_idle <= _mul_6_rshift_idle;
      if(_mul_6_stream_oready) begin
        _mul_6_z_sink_wenable <= 0;
        _mul_6_z_sink_fifo_enq <= 0;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_1 <= _mul_6_stream_ivalid;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_2 <= __mul_6_stream_ivalid_1;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_3 <= __mul_6_stream_ivalid_2;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_4 <= __mul_6_stream_ivalid_3;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_5 <= __mul_6_stream_ivalid_4;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_6 <= __mul_6_stream_ivalid_5;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_7 <= __mul_6_stream_ivalid_6;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_8 <= __mul_6_stream_ivalid_7;
      end 
      if(_mul_6_stream_oready) begin
        _greaterthan_data_125 <= mul_6_rshift_data > 1'sd0;
      end 
      if(_mul_6_stream_oready) begin
        _minus_data_127 <= mul_6_rshift_data - 2'sd1;
      end 
      if(_mul_6_stream_oready) begin
        _greatereq_data_138 <= mul_6_x_data >= 1'sd0;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_696__variable_122 <= mul_6_x_data;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_699__variable_123 <= mul_6_y_data;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_702__variable_124 <= mul_6_rshift_data;
      end 
      if(_mul_6_stream_oready) begin
        _sll_data_129 <= 2'sd1 << _minus_data_127;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_693_greaterthan_125 <= _greaterthan_data_125;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_694_greatereq_138 <= _greatereq_data_138;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_697__delay_696__variable_122 <= __delay_data_696__variable_122;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_700__delay_699__variable_123 <= __delay_data_699__variable_123;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_703__delay_702__variable_124 <= __delay_data_702__variable_124;
      end 
      if(_mul_6_stream_oready) begin
        _cond_data_135 <= (__delay_data_693_greaterthan_125)? _sll_data_129 : 1'sd0;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_695__delay_694_greatereq_138 <= __delay_data_694_greatereq_138;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_698__delay_697__delay_696__variable_122 <= __delay_data_697__delay_696__variable_122;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_701__delay_700__delay_699__variable_123 <= __delay_data_700__delay_699__variable_123;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_704__delay_703__delay_702__variable_124 <= __delay_data_703__delay_702__variable_124;
      end 
      if(_mul_6_stream_oready) begin
        __muladd_madd_odata_reg_141 <= __muladd_madd_odata_141;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_705__delay_704__delay_703____variable_124 <= __delay_data_704__delay_703__delay_702__variable_124;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_706__delay_705__delay_704____variable_124 <= __delay_data_705__delay_704__delay_703____variable_124;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_707__delay_706__delay_705____variable_124 <= __delay_data_706__delay_705__delay_704____variable_124;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_708__delay_707__delay_706____variable_124 <= __delay_data_707__delay_706__delay_705____variable_124;
      end 
      if(_mul_6_stream_oready) begin
        _sra_data_142 <= __muladd_data_141 >>> __delay_data_708__delay_707__delay_706____variable_124;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_122 <= _cond_data_641;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_123 <= __delay_data_960_reinterpretcast_611;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_124 <= _plus_data_709;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_475 <= _mul_6_source_start;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_476 <= _tmp_475;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_477 <= _tmp_476;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_478 <= _mul_6_source_start;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_479 <= _tmp_478;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_480 <= _tmp_479;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_481 <= _tmp_480;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_482 <= _tmp_481;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_483 <= _tmp_482;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_484 <= _tmp_483;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_485 <= _tmp_484;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_486 <= _tmp_485;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_487 <= _tmp_486;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_488 <= _mul_6_source_stop;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_489 <= _tmp_488;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_490 <= _tmp_489;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_491 <= _tmp_490;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_492 <= _tmp_491;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_493 <= _tmp_492;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_494 <= _tmp_493;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_495 <= _tmp_494;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_496 <= _tmp_495;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_497 <= _tmp_496;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_498 <= _mul_6_source_busy;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_499 <= _tmp_498;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_500 <= _tmp_499;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_501 <= _tmp_500;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_502 <= _tmp_501;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_503 <= _tmp_502;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_504 <= _tmp_503;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_505 <= _tmp_504;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_506 <= _tmp_505;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_507 <= _tmp_506;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_508 <= _mul_6_sink_busy;
      end 
      if(!_mul_6_sink_busy && _tmp_508) begin
        _mul_6_busy_reg <= 0;
      end 
      if(_mul_6_source_busy) begin
        _mul_6_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_6_fsm_1 = 1;
  localparam _mul_6_fsm_2 = 2;
  localparam _mul_6_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_6_fsm <= _mul_6_fsm_init;
      _mul_6_source_start <= 0;
      _mul_6_source_busy <= 0;
      _mul_6_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        _mul_6_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_busy) begin
        _mul_6_source_busy <= _stream_conv2d_25_source_busy;
      end 
      if(_mul_6_stream_oready && _tmp_477) begin
        _mul_6_stream_ivalid <= 1;
      end 
      if(_mul_6_stream_oready && 1'd0) begin
        _mul_6_stream_ivalid <= 0;
      end 
      case(_mul_6_fsm)
        _mul_6_fsm_init: begin
          if(_mul_6_run_flag) begin
            _mul_6_source_start <= 1;
          end 
          if(_mul_6_run_flag) begin
            _mul_6_fsm <= _mul_6_fsm_1;
          end 
        end
        _mul_6_fsm_1: begin
          if(_mul_6_source_start && _mul_6_stream_oready) begin
            _mul_6_source_start <= 0;
            _mul_6_source_busy <= 1;
          end 
          if(_mul_6_source_start && _mul_6_stream_oready) begin
            _mul_6_fsm <= _mul_6_fsm_2;
          end 
        end
        _mul_6_fsm_2: begin
          if(_mul_6_stream_oready) begin
            _mul_6_fsm <= _mul_6_fsm_3;
          end 
        end
        _mul_6_fsm_3: begin
          if(_mul_6_stream_oready && 1'd0) begin
            _mul_6_source_busy <= 0;
          end 
          if(_mul_6_stream_oready && 1'd0 && _mul_6_run_flag) begin
            _mul_6_source_start <= 1;
          end 
          if(_mul_6_stream_oready && 1'd0) begin
            _mul_6_fsm <= _mul_6_fsm_init;
          end 
          if(_mul_6_stream_oready && 1'd0 && _mul_6_run_flag) begin
            _mul_6_fsm <= _mul_6_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_7_x_source_ram_renable <= 0;
      _mul_7_x_source_fifo_deq <= 0;
      _mul_7_x_idle <= 1;
      _mul_7_y_source_ram_renable <= 0;
      _mul_7_y_source_fifo_deq <= 0;
      _mul_7_y_idle <= 1;
      _mul_7_rshift_source_ram_renable <= 0;
      _mul_7_rshift_source_fifo_deq <= 0;
      _mul_7_rshift_idle <= 1;
      _mul_7_z_sink_wenable <= 0;
      _mul_7_z_sink_fifo_enq <= 0;
      __mul_7_stream_ivalid_1 <= 0;
      __mul_7_stream_ivalid_2 <= 0;
      __mul_7_stream_ivalid_3 <= 0;
      __mul_7_stream_ivalid_4 <= 0;
      __mul_7_stream_ivalid_5 <= 0;
      __mul_7_stream_ivalid_6 <= 0;
      __mul_7_stream_ivalid_7 <= 0;
      __mul_7_stream_ivalid_8 <= 0;
      _greaterthan_data_146 <= 0;
      _minus_data_148 <= 0;
      _greatereq_data_159 <= 0;
      __delay_data_715__variable_143 <= 0;
      __delay_data_718__variable_144 <= 0;
      __delay_data_721__variable_145 <= 0;
      _sll_data_150 <= 0;
      __delay_data_712_greaterthan_146 <= 0;
      __delay_data_713_greatereq_159 <= 0;
      __delay_data_716__delay_715__variable_143 <= 0;
      __delay_data_719__delay_718__variable_144 <= 0;
      __delay_data_722__delay_721__variable_145 <= 0;
      _cond_data_156 <= 0;
      __delay_data_714__delay_713_greatereq_159 <= 0;
      __delay_data_717__delay_716__delay_715__variable_143 <= 0;
      __delay_data_720__delay_719__delay_718__variable_144 <= 0;
      __delay_data_723__delay_722__delay_721__variable_145 <= 0;
      __muladd_madd_odata_reg_162 <= 0;
      __delay_data_724__delay_723__delay_722____variable_145 <= 0;
      __delay_data_725__delay_724__delay_723____variable_145 <= 0;
      __delay_data_726__delay_725__delay_724____variable_145 <= 0;
      __delay_data_727__delay_726__delay_725____variable_145 <= 0;
      _sra_data_163 <= 0;
      __variable_wdata_143 <= 0;
      __variable_wdata_144 <= 0;
      __variable_wdata_145 <= 0;
      _tmp_509 <= 0;
      _tmp_510 <= 0;
      _tmp_511 <= 0;
      _tmp_512 <= 0;
      _tmp_513 <= 0;
      _tmp_514 <= 0;
      _tmp_515 <= 0;
      _tmp_516 <= 0;
      _tmp_517 <= 0;
      _tmp_518 <= 0;
      _tmp_519 <= 0;
      _tmp_520 <= 0;
      _tmp_521 <= 0;
      _tmp_522 <= 0;
      _tmp_523 <= 0;
      _tmp_524 <= 0;
      _tmp_525 <= 0;
      _tmp_526 <= 0;
      _tmp_527 <= 0;
      _tmp_528 <= 0;
      _tmp_529 <= 0;
      _tmp_530 <= 0;
      _tmp_531 <= 0;
      _tmp_532 <= 0;
      _tmp_533 <= 0;
      _tmp_534 <= 0;
      _tmp_535 <= 0;
      _tmp_536 <= 0;
      _tmp_537 <= 0;
      _tmp_538 <= 0;
      _tmp_539 <= 0;
      _tmp_540 <= 0;
      _tmp_541 <= 0;
      _tmp_542 <= 0;
      _mul_7_busy_reg <= 0;
    end else begin
      if(_mul_7_stream_oready) begin
        _mul_7_x_source_ram_renable <= 0;
        _mul_7_x_source_fifo_deq <= 0;
      end 
      _mul_7_x_idle <= _mul_7_x_idle;
      if(_mul_7_stream_oready) begin
        _mul_7_y_source_ram_renable <= 0;
        _mul_7_y_source_fifo_deq <= 0;
      end 
      _mul_7_y_idle <= _mul_7_y_idle;
      if(_mul_7_stream_oready) begin
        _mul_7_rshift_source_ram_renable <= 0;
        _mul_7_rshift_source_fifo_deq <= 0;
      end 
      _mul_7_rshift_idle <= _mul_7_rshift_idle;
      if(_mul_7_stream_oready) begin
        _mul_7_z_sink_wenable <= 0;
        _mul_7_z_sink_fifo_enq <= 0;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_1 <= _mul_7_stream_ivalid;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_2 <= __mul_7_stream_ivalid_1;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_3 <= __mul_7_stream_ivalid_2;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_4 <= __mul_7_stream_ivalid_3;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_5 <= __mul_7_stream_ivalid_4;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_6 <= __mul_7_stream_ivalid_5;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_7 <= __mul_7_stream_ivalid_6;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_8 <= __mul_7_stream_ivalid_7;
      end 
      if(_mul_7_stream_oready) begin
        _greaterthan_data_146 <= mul_7_rshift_data > 1'sd0;
      end 
      if(_mul_7_stream_oready) begin
        _minus_data_148 <= mul_7_rshift_data - 2'sd1;
      end 
      if(_mul_7_stream_oready) begin
        _greatereq_data_159 <= mul_7_x_data >= 1'sd0;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_715__variable_143 <= mul_7_x_data;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_718__variable_144 <= mul_7_y_data;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_721__variable_145 <= mul_7_rshift_data;
      end 
      if(_mul_7_stream_oready) begin
        _sll_data_150 <= 2'sd1 << _minus_data_148;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_712_greaterthan_146 <= _greaterthan_data_146;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_713_greatereq_159 <= _greatereq_data_159;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_716__delay_715__variable_143 <= __delay_data_715__variable_143;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_719__delay_718__variable_144 <= __delay_data_718__variable_144;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_722__delay_721__variable_145 <= __delay_data_721__variable_145;
      end 
      if(_mul_7_stream_oready) begin
        _cond_data_156 <= (__delay_data_712_greaterthan_146)? _sll_data_150 : 1'sd0;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_714__delay_713_greatereq_159 <= __delay_data_713_greatereq_159;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_717__delay_716__delay_715__variable_143 <= __delay_data_716__delay_715__variable_143;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_720__delay_719__delay_718__variable_144 <= __delay_data_719__delay_718__variable_144;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_723__delay_722__delay_721__variable_145 <= __delay_data_722__delay_721__variable_145;
      end 
      if(_mul_7_stream_oready) begin
        __muladd_madd_odata_reg_162 <= __muladd_madd_odata_162;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_724__delay_723__delay_722____variable_145 <= __delay_data_723__delay_722__delay_721__variable_145;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_725__delay_724__delay_723____variable_145 <= __delay_data_724__delay_723__delay_722____variable_145;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_726__delay_725__delay_724____variable_145 <= __delay_data_725__delay_724__delay_723____variable_145;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_727__delay_726__delay_725____variable_145 <= __delay_data_726__delay_725__delay_724____variable_145;
      end 
      if(_mul_7_stream_oready) begin
        _sra_data_163 <= __muladd_data_162 >>> __delay_data_727__delay_726__delay_725____variable_145;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_143 <= _cond_data_643;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_144 <= __delay_data_962_reinterpretcast_612;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_145 <= _plus_data_728;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_509 <= _mul_7_source_start;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_510 <= _tmp_509;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_511 <= _tmp_510;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_512 <= _mul_7_source_start;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_513 <= _tmp_512;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_514 <= _tmp_513;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_515 <= _tmp_514;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_516 <= _tmp_515;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_517 <= _tmp_516;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_518 <= _tmp_517;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_519 <= _tmp_518;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_520 <= _tmp_519;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_521 <= _tmp_520;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_522 <= _mul_7_source_stop;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_523 <= _tmp_522;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_524 <= _tmp_523;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_525 <= _tmp_524;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_526 <= _tmp_525;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_527 <= _tmp_526;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_528 <= _tmp_527;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_529 <= _tmp_528;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_530 <= _tmp_529;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_531 <= _tmp_530;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_532 <= _mul_7_source_busy;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_533 <= _tmp_532;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_534 <= _tmp_533;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_535 <= _tmp_534;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_536 <= _tmp_535;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_537 <= _tmp_536;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_538 <= _tmp_537;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_539 <= _tmp_538;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_540 <= _tmp_539;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_541 <= _tmp_540;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_542 <= _mul_7_sink_busy;
      end 
      if(!_mul_7_sink_busy && _tmp_542) begin
        _mul_7_busy_reg <= 0;
      end 
      if(_mul_7_source_busy) begin
        _mul_7_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_7_fsm_1 = 1;
  localparam _mul_7_fsm_2 = 2;
  localparam _mul_7_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_7_fsm <= _mul_7_fsm_init;
      _mul_7_source_start <= 0;
      _mul_7_source_busy <= 0;
      _mul_7_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        _mul_7_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_busy) begin
        _mul_7_source_busy <= _stream_conv2d_25_source_busy;
      end 
      if(_mul_7_stream_oready && _tmp_511) begin
        _mul_7_stream_ivalid <= 1;
      end 
      if(_mul_7_stream_oready && 1'd0) begin
        _mul_7_stream_ivalid <= 0;
      end 
      case(_mul_7_fsm)
        _mul_7_fsm_init: begin
          if(_mul_7_run_flag) begin
            _mul_7_source_start <= 1;
          end 
          if(_mul_7_run_flag) begin
            _mul_7_fsm <= _mul_7_fsm_1;
          end 
        end
        _mul_7_fsm_1: begin
          if(_mul_7_source_start && _mul_7_stream_oready) begin
            _mul_7_source_start <= 0;
            _mul_7_source_busy <= 1;
          end 
          if(_mul_7_source_start && _mul_7_stream_oready) begin
            _mul_7_fsm <= _mul_7_fsm_2;
          end 
        end
        _mul_7_fsm_2: begin
          if(_mul_7_stream_oready) begin
            _mul_7_fsm <= _mul_7_fsm_3;
          end 
        end
        _mul_7_fsm_3: begin
          if(_mul_7_stream_oready && 1'd0) begin
            _mul_7_source_busy <= 0;
          end 
          if(_mul_7_stream_oready && 1'd0 && _mul_7_run_flag) begin
            _mul_7_source_start <= 1;
          end 
          if(_mul_7_stream_oready && 1'd0) begin
            _mul_7_fsm <= _mul_7_fsm_init;
          end 
          if(_mul_7_stream_oready && 1'd0 && _mul_7_run_flag) begin
            _mul_7_fsm <= _mul_7_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_8_x_source_ram_renable <= 0;
      _mul_8_x_source_fifo_deq <= 0;
      _mul_8_x_idle <= 1;
      _mul_8_y_source_ram_renable <= 0;
      _mul_8_y_source_fifo_deq <= 0;
      _mul_8_y_idle <= 1;
      _mul_8_rshift_source_ram_renable <= 0;
      _mul_8_rshift_source_fifo_deq <= 0;
      _mul_8_rshift_idle <= 1;
      _mul_8_z_sink_wenable <= 0;
      _mul_8_z_sink_fifo_enq <= 0;
      __mul_8_stream_ivalid_1 <= 0;
      __mul_8_stream_ivalid_2 <= 0;
      __mul_8_stream_ivalid_3 <= 0;
      __mul_8_stream_ivalid_4 <= 0;
      __mul_8_stream_ivalid_5 <= 0;
      __mul_8_stream_ivalid_6 <= 0;
      __mul_8_stream_ivalid_7 <= 0;
      __mul_8_stream_ivalid_8 <= 0;
      _greaterthan_data_167 <= 0;
      _minus_data_169 <= 0;
      _greatereq_data_180 <= 0;
      __delay_data_734__variable_164 <= 0;
      __delay_data_737__variable_165 <= 0;
      __delay_data_740__variable_166 <= 0;
      _sll_data_171 <= 0;
      __delay_data_731_greaterthan_167 <= 0;
      __delay_data_732_greatereq_180 <= 0;
      __delay_data_735__delay_734__variable_164 <= 0;
      __delay_data_738__delay_737__variable_165 <= 0;
      __delay_data_741__delay_740__variable_166 <= 0;
      _cond_data_177 <= 0;
      __delay_data_733__delay_732_greatereq_180 <= 0;
      __delay_data_736__delay_735__delay_734__variable_164 <= 0;
      __delay_data_739__delay_738__delay_737__variable_165 <= 0;
      __delay_data_742__delay_741__delay_740__variable_166 <= 0;
      __muladd_madd_odata_reg_183 <= 0;
      __delay_data_743__delay_742__delay_741____variable_166 <= 0;
      __delay_data_744__delay_743__delay_742____variable_166 <= 0;
      __delay_data_745__delay_744__delay_743____variable_166 <= 0;
      __delay_data_746__delay_745__delay_744____variable_166 <= 0;
      _sra_data_184 <= 0;
      __variable_wdata_164 <= 0;
      __variable_wdata_165 <= 0;
      __variable_wdata_166 <= 0;
      _tmp_543 <= 0;
      _tmp_544 <= 0;
      _tmp_545 <= 0;
      _tmp_546 <= 0;
      _tmp_547 <= 0;
      _tmp_548 <= 0;
      _tmp_549 <= 0;
      _tmp_550 <= 0;
      _tmp_551 <= 0;
      _tmp_552 <= 0;
      _tmp_553 <= 0;
      _tmp_554 <= 0;
      _tmp_555 <= 0;
      _tmp_556 <= 0;
      _tmp_557 <= 0;
      _tmp_558 <= 0;
      _tmp_559 <= 0;
      _tmp_560 <= 0;
      _tmp_561 <= 0;
      _tmp_562 <= 0;
      _tmp_563 <= 0;
      _tmp_564 <= 0;
      _tmp_565 <= 0;
      _tmp_566 <= 0;
      _tmp_567 <= 0;
      _tmp_568 <= 0;
      _tmp_569 <= 0;
      _tmp_570 <= 0;
      _tmp_571 <= 0;
      _tmp_572 <= 0;
      _tmp_573 <= 0;
      _tmp_574 <= 0;
      _tmp_575 <= 0;
      _tmp_576 <= 0;
      _mul_8_busy_reg <= 0;
    end else begin
      if(_mul_8_stream_oready) begin
        _mul_8_x_source_ram_renable <= 0;
        _mul_8_x_source_fifo_deq <= 0;
      end 
      _mul_8_x_idle <= _mul_8_x_idle;
      if(_mul_8_stream_oready) begin
        _mul_8_y_source_ram_renable <= 0;
        _mul_8_y_source_fifo_deq <= 0;
      end 
      _mul_8_y_idle <= _mul_8_y_idle;
      if(_mul_8_stream_oready) begin
        _mul_8_rshift_source_ram_renable <= 0;
        _mul_8_rshift_source_fifo_deq <= 0;
      end 
      _mul_8_rshift_idle <= _mul_8_rshift_idle;
      if(_mul_8_stream_oready) begin
        _mul_8_z_sink_wenable <= 0;
        _mul_8_z_sink_fifo_enq <= 0;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_1 <= _mul_8_stream_ivalid;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_2 <= __mul_8_stream_ivalid_1;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_3 <= __mul_8_stream_ivalid_2;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_4 <= __mul_8_stream_ivalid_3;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_5 <= __mul_8_stream_ivalid_4;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_6 <= __mul_8_stream_ivalid_5;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_7 <= __mul_8_stream_ivalid_6;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_8 <= __mul_8_stream_ivalid_7;
      end 
      if(_mul_8_stream_oready) begin
        _greaterthan_data_167 <= mul_8_rshift_data > 1'sd0;
      end 
      if(_mul_8_stream_oready) begin
        _minus_data_169 <= mul_8_rshift_data - 2'sd1;
      end 
      if(_mul_8_stream_oready) begin
        _greatereq_data_180 <= mul_8_x_data >= 1'sd0;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_734__variable_164 <= mul_8_x_data;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_737__variable_165 <= mul_8_y_data;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_740__variable_166 <= mul_8_rshift_data;
      end 
      if(_mul_8_stream_oready) begin
        _sll_data_171 <= 2'sd1 << _minus_data_169;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_731_greaterthan_167 <= _greaterthan_data_167;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_732_greatereq_180 <= _greatereq_data_180;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_735__delay_734__variable_164 <= __delay_data_734__variable_164;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_738__delay_737__variable_165 <= __delay_data_737__variable_165;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_741__delay_740__variable_166 <= __delay_data_740__variable_166;
      end 
      if(_mul_8_stream_oready) begin
        _cond_data_177 <= (__delay_data_731_greaterthan_167)? _sll_data_171 : 1'sd0;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_733__delay_732_greatereq_180 <= __delay_data_732_greatereq_180;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_736__delay_735__delay_734__variable_164 <= __delay_data_735__delay_734__variable_164;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_739__delay_738__delay_737__variable_165 <= __delay_data_738__delay_737__variable_165;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_742__delay_741__delay_740__variable_166 <= __delay_data_741__delay_740__variable_166;
      end 
      if(_mul_8_stream_oready) begin
        __muladd_madd_odata_reg_183 <= __muladd_madd_odata_183;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_743__delay_742__delay_741____variable_166 <= __delay_data_742__delay_741__delay_740__variable_166;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_744__delay_743__delay_742____variable_166 <= __delay_data_743__delay_742__delay_741____variable_166;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_745__delay_744__delay_743____variable_166 <= __delay_data_744__delay_743__delay_742____variable_166;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_746__delay_745__delay_744____variable_166 <= __delay_data_745__delay_744__delay_743____variable_166;
      end 
      if(_mul_8_stream_oready) begin
        _sra_data_184 <= __muladd_data_183 >>> __delay_data_746__delay_745__delay_744____variable_166;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_164 <= _cond_data_645;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_165 <= __delay_data_964_reinterpretcast_613;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_166 <= _plus_data_747;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_543 <= _mul_8_source_start;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_544 <= _tmp_543;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_545 <= _tmp_544;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_546 <= _mul_8_source_start;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_547 <= _tmp_546;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_548 <= _tmp_547;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_549 <= _tmp_548;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_550 <= _tmp_549;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_551 <= _tmp_550;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_552 <= _tmp_551;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_553 <= _tmp_552;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_554 <= _tmp_553;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_555 <= _tmp_554;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_556 <= _mul_8_source_stop;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_557 <= _tmp_556;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_558 <= _tmp_557;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_559 <= _tmp_558;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_560 <= _tmp_559;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_561 <= _tmp_560;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_562 <= _tmp_561;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_563 <= _tmp_562;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_564 <= _tmp_563;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_565 <= _tmp_564;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_566 <= _mul_8_source_busy;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_567 <= _tmp_566;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_568 <= _tmp_567;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_569 <= _tmp_568;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_570 <= _tmp_569;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_571 <= _tmp_570;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_572 <= _tmp_571;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_573 <= _tmp_572;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_574 <= _tmp_573;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_575 <= _tmp_574;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_576 <= _mul_8_sink_busy;
      end 
      if(!_mul_8_sink_busy && _tmp_576) begin
        _mul_8_busy_reg <= 0;
      end 
      if(_mul_8_source_busy) begin
        _mul_8_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_8_fsm_1 = 1;
  localparam _mul_8_fsm_2 = 2;
  localparam _mul_8_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_8_fsm <= _mul_8_fsm_init;
      _mul_8_source_start <= 0;
      _mul_8_source_busy <= 0;
      _mul_8_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        _mul_8_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_busy) begin
        _mul_8_source_busy <= _stream_conv2d_25_source_busy;
      end 
      if(_mul_8_stream_oready && _tmp_545) begin
        _mul_8_stream_ivalid <= 1;
      end 
      if(_mul_8_stream_oready && 1'd0) begin
        _mul_8_stream_ivalid <= 0;
      end 
      case(_mul_8_fsm)
        _mul_8_fsm_init: begin
          if(_mul_8_run_flag) begin
            _mul_8_source_start <= 1;
          end 
          if(_mul_8_run_flag) begin
            _mul_8_fsm <= _mul_8_fsm_1;
          end 
        end
        _mul_8_fsm_1: begin
          if(_mul_8_source_start && _mul_8_stream_oready) begin
            _mul_8_source_start <= 0;
            _mul_8_source_busy <= 1;
          end 
          if(_mul_8_source_start && _mul_8_stream_oready) begin
            _mul_8_fsm <= _mul_8_fsm_2;
          end 
        end
        _mul_8_fsm_2: begin
          if(_mul_8_stream_oready) begin
            _mul_8_fsm <= _mul_8_fsm_3;
          end 
        end
        _mul_8_fsm_3: begin
          if(_mul_8_stream_oready && 1'd0) begin
            _mul_8_source_busy <= 0;
          end 
          if(_mul_8_stream_oready && 1'd0 && _mul_8_run_flag) begin
            _mul_8_source_start <= 1;
          end 
          if(_mul_8_stream_oready && 1'd0) begin
            _mul_8_fsm <= _mul_8_fsm_init;
          end 
          if(_mul_8_stream_oready && 1'd0 && _mul_8_run_flag) begin
            _mul_8_fsm <= _mul_8_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_9_x_source_ram_renable <= 0;
      _mul_9_x_source_fifo_deq <= 0;
      _mul_9_x_idle <= 1;
      _mul_9_y_source_ram_renable <= 0;
      _mul_9_y_source_fifo_deq <= 0;
      _mul_9_y_idle <= 1;
      _mul_9_rshift_source_ram_renable <= 0;
      _mul_9_rshift_source_fifo_deq <= 0;
      _mul_9_rshift_idle <= 1;
      _mul_9_z_sink_wenable <= 0;
      _mul_9_z_sink_fifo_enq <= 0;
      __mul_9_stream_ivalid_1 <= 0;
      __mul_9_stream_ivalid_2 <= 0;
      __mul_9_stream_ivalid_3 <= 0;
      __mul_9_stream_ivalid_4 <= 0;
      __mul_9_stream_ivalid_5 <= 0;
      __mul_9_stream_ivalid_6 <= 0;
      __mul_9_stream_ivalid_7 <= 0;
      __mul_9_stream_ivalid_8 <= 0;
      _greaterthan_data_188 <= 0;
      _minus_data_190 <= 0;
      _greatereq_data_201 <= 0;
      __delay_data_753__variable_185 <= 0;
      __delay_data_756__variable_186 <= 0;
      __delay_data_759__variable_187 <= 0;
      _sll_data_192 <= 0;
      __delay_data_750_greaterthan_188 <= 0;
      __delay_data_751_greatereq_201 <= 0;
      __delay_data_754__delay_753__variable_185 <= 0;
      __delay_data_757__delay_756__variable_186 <= 0;
      __delay_data_760__delay_759__variable_187 <= 0;
      _cond_data_198 <= 0;
      __delay_data_752__delay_751_greatereq_201 <= 0;
      __delay_data_755__delay_754__delay_753__variable_185 <= 0;
      __delay_data_758__delay_757__delay_756__variable_186 <= 0;
      __delay_data_761__delay_760__delay_759__variable_187 <= 0;
      __muladd_madd_odata_reg_204 <= 0;
      __delay_data_762__delay_761__delay_760____variable_187 <= 0;
      __delay_data_763__delay_762__delay_761____variable_187 <= 0;
      __delay_data_764__delay_763__delay_762____variable_187 <= 0;
      __delay_data_765__delay_764__delay_763____variable_187 <= 0;
      _sra_data_205 <= 0;
      __variable_wdata_185 <= 0;
      __variable_wdata_186 <= 0;
      __variable_wdata_187 <= 0;
      _tmp_577 <= 0;
      _tmp_578 <= 0;
      _tmp_579 <= 0;
      _tmp_580 <= 0;
      _tmp_581 <= 0;
      _tmp_582 <= 0;
      _tmp_583 <= 0;
      _tmp_584 <= 0;
      _tmp_585 <= 0;
      _tmp_586 <= 0;
      _tmp_587 <= 0;
      _tmp_588 <= 0;
      _tmp_589 <= 0;
      _tmp_590 <= 0;
      _tmp_591 <= 0;
      _tmp_592 <= 0;
      _tmp_593 <= 0;
      _tmp_594 <= 0;
      _tmp_595 <= 0;
      _tmp_596 <= 0;
      _tmp_597 <= 0;
      _tmp_598 <= 0;
      _tmp_599 <= 0;
      _tmp_600 <= 0;
      _tmp_601 <= 0;
      _tmp_602 <= 0;
      _tmp_603 <= 0;
      _tmp_604 <= 0;
      _tmp_605 <= 0;
      _tmp_606 <= 0;
      _tmp_607 <= 0;
      _tmp_608 <= 0;
      _tmp_609 <= 0;
      _tmp_610 <= 0;
      _mul_9_busy_reg <= 0;
    end else begin
      if(_mul_9_stream_oready) begin
        _mul_9_x_source_ram_renable <= 0;
        _mul_9_x_source_fifo_deq <= 0;
      end 
      _mul_9_x_idle <= _mul_9_x_idle;
      if(_mul_9_stream_oready) begin
        _mul_9_y_source_ram_renable <= 0;
        _mul_9_y_source_fifo_deq <= 0;
      end 
      _mul_9_y_idle <= _mul_9_y_idle;
      if(_mul_9_stream_oready) begin
        _mul_9_rshift_source_ram_renable <= 0;
        _mul_9_rshift_source_fifo_deq <= 0;
      end 
      _mul_9_rshift_idle <= _mul_9_rshift_idle;
      if(_mul_9_stream_oready) begin
        _mul_9_z_sink_wenable <= 0;
        _mul_9_z_sink_fifo_enq <= 0;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_1 <= _mul_9_stream_ivalid;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_2 <= __mul_9_stream_ivalid_1;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_3 <= __mul_9_stream_ivalid_2;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_4 <= __mul_9_stream_ivalid_3;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_5 <= __mul_9_stream_ivalid_4;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_6 <= __mul_9_stream_ivalid_5;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_7 <= __mul_9_stream_ivalid_6;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_8 <= __mul_9_stream_ivalid_7;
      end 
      if(_mul_9_stream_oready) begin
        _greaterthan_data_188 <= mul_9_rshift_data > 1'sd0;
      end 
      if(_mul_9_stream_oready) begin
        _minus_data_190 <= mul_9_rshift_data - 2'sd1;
      end 
      if(_mul_9_stream_oready) begin
        _greatereq_data_201 <= mul_9_x_data >= 1'sd0;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_753__variable_185 <= mul_9_x_data;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_756__variable_186 <= mul_9_y_data;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_759__variable_187 <= mul_9_rshift_data;
      end 
      if(_mul_9_stream_oready) begin
        _sll_data_192 <= 2'sd1 << _minus_data_190;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_750_greaterthan_188 <= _greaterthan_data_188;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_751_greatereq_201 <= _greatereq_data_201;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_754__delay_753__variable_185 <= __delay_data_753__variable_185;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_757__delay_756__variable_186 <= __delay_data_756__variable_186;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_760__delay_759__variable_187 <= __delay_data_759__variable_187;
      end 
      if(_mul_9_stream_oready) begin
        _cond_data_198 <= (__delay_data_750_greaterthan_188)? _sll_data_192 : 1'sd0;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_752__delay_751_greatereq_201 <= __delay_data_751_greatereq_201;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_755__delay_754__delay_753__variable_185 <= __delay_data_754__delay_753__variable_185;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_758__delay_757__delay_756__variable_186 <= __delay_data_757__delay_756__variable_186;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_761__delay_760__delay_759__variable_187 <= __delay_data_760__delay_759__variable_187;
      end 
      if(_mul_9_stream_oready) begin
        __muladd_madd_odata_reg_204 <= __muladd_madd_odata_204;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_762__delay_761__delay_760____variable_187 <= __delay_data_761__delay_760__delay_759__variable_187;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_763__delay_762__delay_761____variable_187 <= __delay_data_762__delay_761__delay_760____variable_187;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_764__delay_763__delay_762____variable_187 <= __delay_data_763__delay_762__delay_761____variable_187;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_765__delay_764__delay_763____variable_187 <= __delay_data_764__delay_763__delay_762____variable_187;
      end 
      if(_mul_9_stream_oready) begin
        _sra_data_205 <= __muladd_data_204 >>> __delay_data_765__delay_764__delay_763____variable_187;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_185 <= _cond_data_647;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_186 <= __delay_data_966_reinterpretcast_614;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_187 <= _plus_data_766;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_577 <= _mul_9_source_start;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_578 <= _tmp_577;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_579 <= _tmp_578;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_580 <= _mul_9_source_start;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_581 <= _tmp_580;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_582 <= _tmp_581;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_583 <= _tmp_582;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_584 <= _tmp_583;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_585 <= _tmp_584;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_586 <= _tmp_585;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_587 <= _tmp_586;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_588 <= _tmp_587;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_589 <= _tmp_588;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_590 <= _mul_9_source_stop;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_591 <= _tmp_590;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_592 <= _tmp_591;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_593 <= _tmp_592;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_594 <= _tmp_593;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_595 <= _tmp_594;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_596 <= _tmp_595;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_597 <= _tmp_596;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_598 <= _tmp_597;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_599 <= _tmp_598;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_600 <= _mul_9_source_busy;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_601 <= _tmp_600;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_602 <= _tmp_601;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_603 <= _tmp_602;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_604 <= _tmp_603;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_605 <= _tmp_604;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_606 <= _tmp_605;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_607 <= _tmp_606;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_608 <= _tmp_607;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_609 <= _tmp_608;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_610 <= _mul_9_sink_busy;
      end 
      if(!_mul_9_sink_busy && _tmp_610) begin
        _mul_9_busy_reg <= 0;
      end 
      if(_mul_9_source_busy) begin
        _mul_9_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_9_fsm_1 = 1;
  localparam _mul_9_fsm_2 = 2;
  localparam _mul_9_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_9_fsm <= _mul_9_fsm_init;
      _mul_9_source_start <= 0;
      _mul_9_source_busy <= 0;
      _mul_9_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        _mul_9_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_busy) begin
        _mul_9_source_busy <= _stream_conv2d_25_source_busy;
      end 
      if(_mul_9_stream_oready && _tmp_579) begin
        _mul_9_stream_ivalid <= 1;
      end 
      if(_mul_9_stream_oready && 1'd0) begin
        _mul_9_stream_ivalid <= 0;
      end 
      case(_mul_9_fsm)
        _mul_9_fsm_init: begin
          if(_mul_9_run_flag) begin
            _mul_9_source_start <= 1;
          end 
          if(_mul_9_run_flag) begin
            _mul_9_fsm <= _mul_9_fsm_1;
          end 
        end
        _mul_9_fsm_1: begin
          if(_mul_9_source_start && _mul_9_stream_oready) begin
            _mul_9_source_start <= 0;
            _mul_9_source_busy <= 1;
          end 
          if(_mul_9_source_start && _mul_9_stream_oready) begin
            _mul_9_fsm <= _mul_9_fsm_2;
          end 
        end
        _mul_9_fsm_2: begin
          if(_mul_9_stream_oready) begin
            _mul_9_fsm <= _mul_9_fsm_3;
          end 
        end
        _mul_9_fsm_3: begin
          if(_mul_9_stream_oready && 1'd0) begin
            _mul_9_source_busy <= 0;
          end 
          if(_mul_9_stream_oready && 1'd0 && _mul_9_run_flag) begin
            _mul_9_source_start <= 1;
          end 
          if(_mul_9_stream_oready && 1'd0) begin
            _mul_9_fsm <= _mul_9_fsm_init;
          end 
          if(_mul_9_stream_oready && 1'd0 && _mul_9_run_flag) begin
            _mul_9_fsm <= _mul_9_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_10_x_source_ram_renable <= 0;
      _mul_10_x_source_fifo_deq <= 0;
      _mul_10_x_idle <= 1;
      _mul_10_y_source_ram_renable <= 0;
      _mul_10_y_source_fifo_deq <= 0;
      _mul_10_y_idle <= 1;
      _mul_10_rshift_source_ram_renable <= 0;
      _mul_10_rshift_source_fifo_deq <= 0;
      _mul_10_rshift_idle <= 1;
      _mul_10_z_sink_wenable <= 0;
      _mul_10_z_sink_fifo_enq <= 0;
      __mul_10_stream_ivalid_1 <= 0;
      __mul_10_stream_ivalid_2 <= 0;
      __mul_10_stream_ivalid_3 <= 0;
      __mul_10_stream_ivalid_4 <= 0;
      __mul_10_stream_ivalid_5 <= 0;
      __mul_10_stream_ivalid_6 <= 0;
      __mul_10_stream_ivalid_7 <= 0;
      __mul_10_stream_ivalid_8 <= 0;
      _greaterthan_data_209 <= 0;
      _minus_data_211 <= 0;
      _greatereq_data_222 <= 0;
      __delay_data_772__variable_206 <= 0;
      __delay_data_775__variable_207 <= 0;
      __delay_data_778__variable_208 <= 0;
      _sll_data_213 <= 0;
      __delay_data_769_greaterthan_209 <= 0;
      __delay_data_770_greatereq_222 <= 0;
      __delay_data_773__delay_772__variable_206 <= 0;
      __delay_data_776__delay_775__variable_207 <= 0;
      __delay_data_779__delay_778__variable_208 <= 0;
      _cond_data_219 <= 0;
      __delay_data_771__delay_770_greatereq_222 <= 0;
      __delay_data_774__delay_773__delay_772__variable_206 <= 0;
      __delay_data_777__delay_776__delay_775__variable_207 <= 0;
      __delay_data_780__delay_779__delay_778__variable_208 <= 0;
      __muladd_madd_odata_reg_225 <= 0;
      __delay_data_781__delay_780__delay_779____variable_208 <= 0;
      __delay_data_782__delay_781__delay_780____variable_208 <= 0;
      __delay_data_783__delay_782__delay_781____variable_208 <= 0;
      __delay_data_784__delay_783__delay_782____variable_208 <= 0;
      _sra_data_226 <= 0;
      __variable_wdata_206 <= 0;
      __variable_wdata_207 <= 0;
      __variable_wdata_208 <= 0;
      _tmp_611 <= 0;
      _tmp_612 <= 0;
      _tmp_613 <= 0;
      _tmp_614 <= 0;
      _tmp_615 <= 0;
      _tmp_616 <= 0;
      _tmp_617 <= 0;
      _tmp_618 <= 0;
      _tmp_619 <= 0;
      _tmp_620 <= 0;
      _tmp_621 <= 0;
      _tmp_622 <= 0;
      _tmp_623 <= 0;
      _tmp_624 <= 0;
      _tmp_625 <= 0;
      _tmp_626 <= 0;
      _tmp_627 <= 0;
      _tmp_628 <= 0;
      _tmp_629 <= 0;
      _tmp_630 <= 0;
      _tmp_631 <= 0;
      _tmp_632 <= 0;
      _tmp_633 <= 0;
      _tmp_634 <= 0;
      _tmp_635 <= 0;
      _tmp_636 <= 0;
      _tmp_637 <= 0;
      _tmp_638 <= 0;
      _tmp_639 <= 0;
      _tmp_640 <= 0;
      _tmp_641 <= 0;
      _tmp_642 <= 0;
      _tmp_643 <= 0;
      _tmp_644 <= 0;
      _mul_10_busy_reg <= 0;
    end else begin
      if(_mul_10_stream_oready) begin
        _mul_10_x_source_ram_renable <= 0;
        _mul_10_x_source_fifo_deq <= 0;
      end 
      _mul_10_x_idle <= _mul_10_x_idle;
      if(_mul_10_stream_oready) begin
        _mul_10_y_source_ram_renable <= 0;
        _mul_10_y_source_fifo_deq <= 0;
      end 
      _mul_10_y_idle <= _mul_10_y_idle;
      if(_mul_10_stream_oready) begin
        _mul_10_rshift_source_ram_renable <= 0;
        _mul_10_rshift_source_fifo_deq <= 0;
      end 
      _mul_10_rshift_idle <= _mul_10_rshift_idle;
      if(_mul_10_stream_oready) begin
        _mul_10_z_sink_wenable <= 0;
        _mul_10_z_sink_fifo_enq <= 0;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_1 <= _mul_10_stream_ivalid;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_2 <= __mul_10_stream_ivalid_1;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_3 <= __mul_10_stream_ivalid_2;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_4 <= __mul_10_stream_ivalid_3;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_5 <= __mul_10_stream_ivalid_4;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_6 <= __mul_10_stream_ivalid_5;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_7 <= __mul_10_stream_ivalid_6;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_8 <= __mul_10_stream_ivalid_7;
      end 
      if(_mul_10_stream_oready) begin
        _greaterthan_data_209 <= mul_10_rshift_data > 1'sd0;
      end 
      if(_mul_10_stream_oready) begin
        _minus_data_211 <= mul_10_rshift_data - 2'sd1;
      end 
      if(_mul_10_stream_oready) begin
        _greatereq_data_222 <= mul_10_x_data >= 1'sd0;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_772__variable_206 <= mul_10_x_data;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_775__variable_207 <= mul_10_y_data;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_778__variable_208 <= mul_10_rshift_data;
      end 
      if(_mul_10_stream_oready) begin
        _sll_data_213 <= 2'sd1 << _minus_data_211;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_769_greaterthan_209 <= _greaterthan_data_209;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_770_greatereq_222 <= _greatereq_data_222;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_773__delay_772__variable_206 <= __delay_data_772__variable_206;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_776__delay_775__variable_207 <= __delay_data_775__variable_207;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_779__delay_778__variable_208 <= __delay_data_778__variable_208;
      end 
      if(_mul_10_stream_oready) begin
        _cond_data_219 <= (__delay_data_769_greaterthan_209)? _sll_data_213 : 1'sd0;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_771__delay_770_greatereq_222 <= __delay_data_770_greatereq_222;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_774__delay_773__delay_772__variable_206 <= __delay_data_773__delay_772__variable_206;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_777__delay_776__delay_775__variable_207 <= __delay_data_776__delay_775__variable_207;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_780__delay_779__delay_778__variable_208 <= __delay_data_779__delay_778__variable_208;
      end 
      if(_mul_10_stream_oready) begin
        __muladd_madd_odata_reg_225 <= __muladd_madd_odata_225;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_781__delay_780__delay_779____variable_208 <= __delay_data_780__delay_779__delay_778__variable_208;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_782__delay_781__delay_780____variable_208 <= __delay_data_781__delay_780__delay_779____variable_208;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_783__delay_782__delay_781____variable_208 <= __delay_data_782__delay_781__delay_780____variable_208;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_784__delay_783__delay_782____variable_208 <= __delay_data_783__delay_782__delay_781____variable_208;
      end 
      if(_mul_10_stream_oready) begin
        _sra_data_226 <= __muladd_data_225 >>> __delay_data_784__delay_783__delay_782____variable_208;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_206 <= _cond_data_649;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_207 <= __delay_data_968_reinterpretcast_615;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_208 <= _plus_data_785;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_611 <= _mul_10_source_start;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_612 <= _tmp_611;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_613 <= _tmp_612;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_614 <= _mul_10_source_start;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_615 <= _tmp_614;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_616 <= _tmp_615;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_617 <= _tmp_616;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_618 <= _tmp_617;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_619 <= _tmp_618;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_620 <= _tmp_619;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_621 <= _tmp_620;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_622 <= _tmp_621;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_623 <= _tmp_622;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_624 <= _mul_10_source_stop;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_625 <= _tmp_624;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_626 <= _tmp_625;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_627 <= _tmp_626;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_628 <= _tmp_627;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_629 <= _tmp_628;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_630 <= _tmp_629;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_631 <= _tmp_630;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_632 <= _tmp_631;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_633 <= _tmp_632;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_634 <= _mul_10_source_busy;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_635 <= _tmp_634;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_636 <= _tmp_635;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_637 <= _tmp_636;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_638 <= _tmp_637;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_639 <= _tmp_638;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_640 <= _tmp_639;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_641 <= _tmp_640;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_642 <= _tmp_641;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_643 <= _tmp_642;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_644 <= _mul_10_sink_busy;
      end 
      if(!_mul_10_sink_busy && _tmp_644) begin
        _mul_10_busy_reg <= 0;
      end 
      if(_mul_10_source_busy) begin
        _mul_10_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_10_fsm_1 = 1;
  localparam _mul_10_fsm_2 = 2;
  localparam _mul_10_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_10_fsm <= _mul_10_fsm_init;
      _mul_10_source_start <= 0;
      _mul_10_source_busy <= 0;
      _mul_10_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        _mul_10_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_busy) begin
        _mul_10_source_busy <= _stream_conv2d_25_source_busy;
      end 
      if(_mul_10_stream_oready && _tmp_613) begin
        _mul_10_stream_ivalid <= 1;
      end 
      if(_mul_10_stream_oready && 1'd0) begin
        _mul_10_stream_ivalid <= 0;
      end 
      case(_mul_10_fsm)
        _mul_10_fsm_init: begin
          if(_mul_10_run_flag) begin
            _mul_10_source_start <= 1;
          end 
          if(_mul_10_run_flag) begin
            _mul_10_fsm <= _mul_10_fsm_1;
          end 
        end
        _mul_10_fsm_1: begin
          if(_mul_10_source_start && _mul_10_stream_oready) begin
            _mul_10_source_start <= 0;
            _mul_10_source_busy <= 1;
          end 
          if(_mul_10_source_start && _mul_10_stream_oready) begin
            _mul_10_fsm <= _mul_10_fsm_2;
          end 
        end
        _mul_10_fsm_2: begin
          if(_mul_10_stream_oready) begin
            _mul_10_fsm <= _mul_10_fsm_3;
          end 
        end
        _mul_10_fsm_3: begin
          if(_mul_10_stream_oready && 1'd0) begin
            _mul_10_source_busy <= 0;
          end 
          if(_mul_10_stream_oready && 1'd0 && _mul_10_run_flag) begin
            _mul_10_source_start <= 1;
          end 
          if(_mul_10_stream_oready && 1'd0) begin
            _mul_10_fsm <= _mul_10_fsm_init;
          end 
          if(_mul_10_stream_oready && 1'd0 && _mul_10_run_flag) begin
            _mul_10_fsm <= _mul_10_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_11_x_source_ram_renable <= 0;
      _mul_11_x_source_fifo_deq <= 0;
      _mul_11_x_idle <= 1;
      _mul_11_y_source_ram_renable <= 0;
      _mul_11_y_source_fifo_deq <= 0;
      _mul_11_y_idle <= 1;
      _mul_11_rshift_source_ram_renable <= 0;
      _mul_11_rshift_source_fifo_deq <= 0;
      _mul_11_rshift_idle <= 1;
      _mul_11_z_sink_wenable <= 0;
      _mul_11_z_sink_fifo_enq <= 0;
      __mul_11_stream_ivalid_1 <= 0;
      __mul_11_stream_ivalid_2 <= 0;
      __mul_11_stream_ivalid_3 <= 0;
      __mul_11_stream_ivalid_4 <= 0;
      __mul_11_stream_ivalid_5 <= 0;
      __mul_11_stream_ivalid_6 <= 0;
      __mul_11_stream_ivalid_7 <= 0;
      __mul_11_stream_ivalid_8 <= 0;
      _greaterthan_data_230 <= 0;
      _minus_data_232 <= 0;
      _greatereq_data_243 <= 0;
      __delay_data_791__variable_227 <= 0;
      __delay_data_794__variable_228 <= 0;
      __delay_data_797__variable_229 <= 0;
      _sll_data_234 <= 0;
      __delay_data_788_greaterthan_230 <= 0;
      __delay_data_789_greatereq_243 <= 0;
      __delay_data_792__delay_791__variable_227 <= 0;
      __delay_data_795__delay_794__variable_228 <= 0;
      __delay_data_798__delay_797__variable_229 <= 0;
      _cond_data_240 <= 0;
      __delay_data_790__delay_789_greatereq_243 <= 0;
      __delay_data_793__delay_792__delay_791__variable_227 <= 0;
      __delay_data_796__delay_795__delay_794__variable_228 <= 0;
      __delay_data_799__delay_798__delay_797__variable_229 <= 0;
      __muladd_madd_odata_reg_246 <= 0;
      __delay_data_800__delay_799__delay_798____variable_229 <= 0;
      __delay_data_801__delay_800__delay_799____variable_229 <= 0;
      __delay_data_802__delay_801__delay_800____variable_229 <= 0;
      __delay_data_803__delay_802__delay_801____variable_229 <= 0;
      _sra_data_247 <= 0;
      __variable_wdata_227 <= 0;
      __variable_wdata_228 <= 0;
      __variable_wdata_229 <= 0;
      _tmp_645 <= 0;
      _tmp_646 <= 0;
      _tmp_647 <= 0;
      _tmp_648 <= 0;
      _tmp_649 <= 0;
      _tmp_650 <= 0;
      _tmp_651 <= 0;
      _tmp_652 <= 0;
      _tmp_653 <= 0;
      _tmp_654 <= 0;
      _tmp_655 <= 0;
      _tmp_656 <= 0;
      _tmp_657 <= 0;
      _tmp_658 <= 0;
      _tmp_659 <= 0;
      _tmp_660 <= 0;
      _tmp_661 <= 0;
      _tmp_662 <= 0;
      _tmp_663 <= 0;
      _tmp_664 <= 0;
      _tmp_665 <= 0;
      _tmp_666 <= 0;
      _tmp_667 <= 0;
      _tmp_668 <= 0;
      _tmp_669 <= 0;
      _tmp_670 <= 0;
      _tmp_671 <= 0;
      _tmp_672 <= 0;
      _tmp_673 <= 0;
      _tmp_674 <= 0;
      _tmp_675 <= 0;
      _tmp_676 <= 0;
      _tmp_677 <= 0;
      _tmp_678 <= 0;
      _mul_11_busy_reg <= 0;
    end else begin
      if(_mul_11_stream_oready) begin
        _mul_11_x_source_ram_renable <= 0;
        _mul_11_x_source_fifo_deq <= 0;
      end 
      _mul_11_x_idle <= _mul_11_x_idle;
      if(_mul_11_stream_oready) begin
        _mul_11_y_source_ram_renable <= 0;
        _mul_11_y_source_fifo_deq <= 0;
      end 
      _mul_11_y_idle <= _mul_11_y_idle;
      if(_mul_11_stream_oready) begin
        _mul_11_rshift_source_ram_renable <= 0;
        _mul_11_rshift_source_fifo_deq <= 0;
      end 
      _mul_11_rshift_idle <= _mul_11_rshift_idle;
      if(_mul_11_stream_oready) begin
        _mul_11_z_sink_wenable <= 0;
        _mul_11_z_sink_fifo_enq <= 0;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_1 <= _mul_11_stream_ivalid;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_2 <= __mul_11_stream_ivalid_1;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_3 <= __mul_11_stream_ivalid_2;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_4 <= __mul_11_stream_ivalid_3;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_5 <= __mul_11_stream_ivalid_4;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_6 <= __mul_11_stream_ivalid_5;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_7 <= __mul_11_stream_ivalid_6;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_8 <= __mul_11_stream_ivalid_7;
      end 
      if(_mul_11_stream_oready) begin
        _greaterthan_data_230 <= mul_11_rshift_data > 1'sd0;
      end 
      if(_mul_11_stream_oready) begin
        _minus_data_232 <= mul_11_rshift_data - 2'sd1;
      end 
      if(_mul_11_stream_oready) begin
        _greatereq_data_243 <= mul_11_x_data >= 1'sd0;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_791__variable_227 <= mul_11_x_data;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_794__variable_228 <= mul_11_y_data;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_797__variable_229 <= mul_11_rshift_data;
      end 
      if(_mul_11_stream_oready) begin
        _sll_data_234 <= 2'sd1 << _minus_data_232;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_788_greaterthan_230 <= _greaterthan_data_230;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_789_greatereq_243 <= _greatereq_data_243;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_792__delay_791__variable_227 <= __delay_data_791__variable_227;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_795__delay_794__variable_228 <= __delay_data_794__variable_228;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_798__delay_797__variable_229 <= __delay_data_797__variable_229;
      end 
      if(_mul_11_stream_oready) begin
        _cond_data_240 <= (__delay_data_788_greaterthan_230)? _sll_data_234 : 1'sd0;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_790__delay_789_greatereq_243 <= __delay_data_789_greatereq_243;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_793__delay_792__delay_791__variable_227 <= __delay_data_792__delay_791__variable_227;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_796__delay_795__delay_794__variable_228 <= __delay_data_795__delay_794__variable_228;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_799__delay_798__delay_797__variable_229 <= __delay_data_798__delay_797__variable_229;
      end 
      if(_mul_11_stream_oready) begin
        __muladd_madd_odata_reg_246 <= __muladd_madd_odata_246;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_800__delay_799__delay_798____variable_229 <= __delay_data_799__delay_798__delay_797__variable_229;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_801__delay_800__delay_799____variable_229 <= __delay_data_800__delay_799__delay_798____variable_229;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_802__delay_801__delay_800____variable_229 <= __delay_data_801__delay_800__delay_799____variable_229;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_803__delay_802__delay_801____variable_229 <= __delay_data_802__delay_801__delay_800____variable_229;
      end 
      if(_mul_11_stream_oready) begin
        _sra_data_247 <= __muladd_data_246 >>> __delay_data_803__delay_802__delay_801____variable_229;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_227 <= _cond_data_651;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_228 <= __delay_data_970_reinterpretcast_616;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_229 <= _plus_data_804;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_645 <= _mul_11_source_start;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_646 <= _tmp_645;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_647 <= _tmp_646;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_648 <= _mul_11_source_start;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_649 <= _tmp_648;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_650 <= _tmp_649;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_651 <= _tmp_650;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_652 <= _tmp_651;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_653 <= _tmp_652;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_654 <= _tmp_653;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_655 <= _tmp_654;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_656 <= _tmp_655;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_657 <= _tmp_656;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_658 <= _mul_11_source_stop;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_659 <= _tmp_658;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_660 <= _tmp_659;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_661 <= _tmp_660;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_662 <= _tmp_661;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_663 <= _tmp_662;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_664 <= _tmp_663;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_665 <= _tmp_664;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_666 <= _tmp_665;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_667 <= _tmp_666;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_668 <= _mul_11_source_busy;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_669 <= _tmp_668;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_670 <= _tmp_669;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_671 <= _tmp_670;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_672 <= _tmp_671;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_673 <= _tmp_672;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_674 <= _tmp_673;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_675 <= _tmp_674;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_676 <= _tmp_675;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_677 <= _tmp_676;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_678 <= _mul_11_sink_busy;
      end 
      if(!_mul_11_sink_busy && _tmp_678) begin
        _mul_11_busy_reg <= 0;
      end 
      if(_mul_11_source_busy) begin
        _mul_11_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_11_fsm_1 = 1;
  localparam _mul_11_fsm_2 = 2;
  localparam _mul_11_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_11_fsm <= _mul_11_fsm_init;
      _mul_11_source_start <= 0;
      _mul_11_source_busy <= 0;
      _mul_11_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        _mul_11_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_busy) begin
        _mul_11_source_busy <= _stream_conv2d_25_source_busy;
      end 
      if(_mul_11_stream_oready && _tmp_647) begin
        _mul_11_stream_ivalid <= 1;
      end 
      if(_mul_11_stream_oready && 1'd0) begin
        _mul_11_stream_ivalid <= 0;
      end 
      case(_mul_11_fsm)
        _mul_11_fsm_init: begin
          if(_mul_11_run_flag) begin
            _mul_11_source_start <= 1;
          end 
          if(_mul_11_run_flag) begin
            _mul_11_fsm <= _mul_11_fsm_1;
          end 
        end
        _mul_11_fsm_1: begin
          if(_mul_11_source_start && _mul_11_stream_oready) begin
            _mul_11_source_start <= 0;
            _mul_11_source_busy <= 1;
          end 
          if(_mul_11_source_start && _mul_11_stream_oready) begin
            _mul_11_fsm <= _mul_11_fsm_2;
          end 
        end
        _mul_11_fsm_2: begin
          if(_mul_11_stream_oready) begin
            _mul_11_fsm <= _mul_11_fsm_3;
          end 
        end
        _mul_11_fsm_3: begin
          if(_mul_11_stream_oready && 1'd0) begin
            _mul_11_source_busy <= 0;
          end 
          if(_mul_11_stream_oready && 1'd0 && _mul_11_run_flag) begin
            _mul_11_source_start <= 1;
          end 
          if(_mul_11_stream_oready && 1'd0) begin
            _mul_11_fsm <= _mul_11_fsm_init;
          end 
          if(_mul_11_stream_oready && 1'd0 && _mul_11_run_flag) begin
            _mul_11_fsm <= _mul_11_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_12_x_source_ram_renable <= 0;
      _mul_12_x_source_fifo_deq <= 0;
      _mul_12_x_idle <= 1;
      _mul_12_y_source_ram_renable <= 0;
      _mul_12_y_source_fifo_deq <= 0;
      _mul_12_y_idle <= 1;
      _mul_12_rshift_source_ram_renable <= 0;
      _mul_12_rshift_source_fifo_deq <= 0;
      _mul_12_rshift_idle <= 1;
      _mul_12_z_sink_wenable <= 0;
      _mul_12_z_sink_fifo_enq <= 0;
      __mul_12_stream_ivalid_1 <= 0;
      __mul_12_stream_ivalid_2 <= 0;
      __mul_12_stream_ivalid_3 <= 0;
      __mul_12_stream_ivalid_4 <= 0;
      __mul_12_stream_ivalid_5 <= 0;
      __mul_12_stream_ivalid_6 <= 0;
      __mul_12_stream_ivalid_7 <= 0;
      __mul_12_stream_ivalid_8 <= 0;
      _greaterthan_data_251 <= 0;
      _minus_data_253 <= 0;
      _greatereq_data_264 <= 0;
      __delay_data_810__variable_248 <= 0;
      __delay_data_813__variable_249 <= 0;
      __delay_data_816__variable_250 <= 0;
      _sll_data_255 <= 0;
      __delay_data_807_greaterthan_251 <= 0;
      __delay_data_808_greatereq_264 <= 0;
      __delay_data_811__delay_810__variable_248 <= 0;
      __delay_data_814__delay_813__variable_249 <= 0;
      __delay_data_817__delay_816__variable_250 <= 0;
      _cond_data_261 <= 0;
      __delay_data_809__delay_808_greatereq_264 <= 0;
      __delay_data_812__delay_811__delay_810__variable_248 <= 0;
      __delay_data_815__delay_814__delay_813__variable_249 <= 0;
      __delay_data_818__delay_817__delay_816__variable_250 <= 0;
      __muladd_madd_odata_reg_267 <= 0;
      __delay_data_819__delay_818__delay_817____variable_250 <= 0;
      __delay_data_820__delay_819__delay_818____variable_250 <= 0;
      __delay_data_821__delay_820__delay_819____variable_250 <= 0;
      __delay_data_822__delay_821__delay_820____variable_250 <= 0;
      _sra_data_268 <= 0;
      __variable_wdata_248 <= 0;
      __variable_wdata_249 <= 0;
      __variable_wdata_250 <= 0;
      _tmp_679 <= 0;
      _tmp_680 <= 0;
      _tmp_681 <= 0;
      _tmp_682 <= 0;
      _tmp_683 <= 0;
      _tmp_684 <= 0;
      _tmp_685 <= 0;
      _tmp_686 <= 0;
      _tmp_687 <= 0;
      _tmp_688 <= 0;
      _tmp_689 <= 0;
      _tmp_690 <= 0;
      _tmp_691 <= 0;
      _tmp_692 <= 0;
      _tmp_693 <= 0;
      _tmp_694 <= 0;
      _tmp_695 <= 0;
      _tmp_696 <= 0;
      _tmp_697 <= 0;
      _tmp_698 <= 0;
      _tmp_699 <= 0;
      _tmp_700 <= 0;
      _tmp_701 <= 0;
      _tmp_702 <= 0;
      _tmp_703 <= 0;
      _tmp_704 <= 0;
      _tmp_705 <= 0;
      _tmp_706 <= 0;
      _tmp_707 <= 0;
      _tmp_708 <= 0;
      _tmp_709 <= 0;
      _tmp_710 <= 0;
      _tmp_711 <= 0;
      _tmp_712 <= 0;
      _mul_12_busy_reg <= 0;
    end else begin
      if(_mul_12_stream_oready) begin
        _mul_12_x_source_ram_renable <= 0;
        _mul_12_x_source_fifo_deq <= 0;
      end 
      _mul_12_x_idle <= _mul_12_x_idle;
      if(_mul_12_stream_oready) begin
        _mul_12_y_source_ram_renable <= 0;
        _mul_12_y_source_fifo_deq <= 0;
      end 
      _mul_12_y_idle <= _mul_12_y_idle;
      if(_mul_12_stream_oready) begin
        _mul_12_rshift_source_ram_renable <= 0;
        _mul_12_rshift_source_fifo_deq <= 0;
      end 
      _mul_12_rshift_idle <= _mul_12_rshift_idle;
      if(_mul_12_stream_oready) begin
        _mul_12_z_sink_wenable <= 0;
        _mul_12_z_sink_fifo_enq <= 0;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_1 <= _mul_12_stream_ivalid;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_2 <= __mul_12_stream_ivalid_1;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_3 <= __mul_12_stream_ivalid_2;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_4 <= __mul_12_stream_ivalid_3;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_5 <= __mul_12_stream_ivalid_4;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_6 <= __mul_12_stream_ivalid_5;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_7 <= __mul_12_stream_ivalid_6;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_8 <= __mul_12_stream_ivalid_7;
      end 
      if(_mul_12_stream_oready) begin
        _greaterthan_data_251 <= mul_12_rshift_data > 1'sd0;
      end 
      if(_mul_12_stream_oready) begin
        _minus_data_253 <= mul_12_rshift_data - 2'sd1;
      end 
      if(_mul_12_stream_oready) begin
        _greatereq_data_264 <= mul_12_x_data >= 1'sd0;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_810__variable_248 <= mul_12_x_data;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_813__variable_249 <= mul_12_y_data;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_816__variable_250 <= mul_12_rshift_data;
      end 
      if(_mul_12_stream_oready) begin
        _sll_data_255 <= 2'sd1 << _minus_data_253;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_807_greaterthan_251 <= _greaterthan_data_251;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_808_greatereq_264 <= _greatereq_data_264;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_811__delay_810__variable_248 <= __delay_data_810__variable_248;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_814__delay_813__variable_249 <= __delay_data_813__variable_249;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_817__delay_816__variable_250 <= __delay_data_816__variable_250;
      end 
      if(_mul_12_stream_oready) begin
        _cond_data_261 <= (__delay_data_807_greaterthan_251)? _sll_data_255 : 1'sd0;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_809__delay_808_greatereq_264 <= __delay_data_808_greatereq_264;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_812__delay_811__delay_810__variable_248 <= __delay_data_811__delay_810__variable_248;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_815__delay_814__delay_813__variable_249 <= __delay_data_814__delay_813__variable_249;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_818__delay_817__delay_816__variable_250 <= __delay_data_817__delay_816__variable_250;
      end 
      if(_mul_12_stream_oready) begin
        __muladd_madd_odata_reg_267 <= __muladd_madd_odata_267;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_819__delay_818__delay_817____variable_250 <= __delay_data_818__delay_817__delay_816__variable_250;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_820__delay_819__delay_818____variable_250 <= __delay_data_819__delay_818__delay_817____variable_250;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_821__delay_820__delay_819____variable_250 <= __delay_data_820__delay_819__delay_818____variable_250;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_822__delay_821__delay_820____variable_250 <= __delay_data_821__delay_820__delay_819____variable_250;
      end 
      if(_mul_12_stream_oready) begin
        _sra_data_268 <= __muladd_data_267 >>> __delay_data_822__delay_821__delay_820____variable_250;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_248 <= _cond_data_653;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_249 <= __delay_data_972_reinterpretcast_617;
      end 
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        __variable_wdata_250 <= _plus_data_823;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_679 <= _mul_12_source_start;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_680 <= _tmp_679;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_681 <= _tmp_680;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_682 <= _mul_12_source_start;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_683 <= _tmp_682;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_684 <= _tmp_683;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_685 <= _tmp_684;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_686 <= _tmp_685;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_687 <= _tmp_686;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_688 <= _tmp_687;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_689 <= _tmp_688;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_690 <= _tmp_689;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_691 <= _tmp_690;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_692 <= _mul_12_source_stop;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_693 <= _tmp_692;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_694 <= _tmp_693;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_695 <= _tmp_694;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_696 <= _tmp_695;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_697 <= _tmp_696;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_698 <= _tmp_697;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_699 <= _tmp_698;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_700 <= _tmp_699;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_701 <= _tmp_700;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_702 <= _mul_12_source_busy;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_703 <= _tmp_702;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_704 <= _tmp_703;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_705 <= _tmp_704;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_706 <= _tmp_705;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_707 <= _tmp_706;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_708 <= _tmp_707;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_709 <= _tmp_708;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_710 <= _tmp_709;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_711 <= _tmp_710;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_712 <= _mul_12_sink_busy;
      end 
      if(!_mul_12_sink_busy && _tmp_712) begin
        _mul_12_busy_reg <= 0;
      end 
      if(_mul_12_source_busy) begin
        _mul_12_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_12_fsm_1 = 1;
  localparam _mul_12_fsm_2 = 2;
  localparam _mul_12_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_12_fsm <= _mul_12_fsm_init;
      _mul_12_source_start <= 0;
      _mul_12_source_busy <= 0;
      _mul_12_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_25_stream_ivalid_1 && _stream_conv2d_25_stream_oready) begin
        _mul_12_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_busy) begin
        _mul_12_source_busy <= _stream_conv2d_25_source_busy;
      end 
      if(_mul_12_stream_oready && _tmp_681) begin
        _mul_12_stream_ivalid <= 1;
      end 
      if(_mul_12_stream_oready && 1'd0) begin
        _mul_12_stream_ivalid <= 0;
      end 
      case(_mul_12_fsm)
        _mul_12_fsm_init: begin
          if(_mul_12_run_flag) begin
            _mul_12_source_start <= 1;
          end 
          if(_mul_12_run_flag) begin
            _mul_12_fsm <= _mul_12_fsm_1;
          end 
        end
        _mul_12_fsm_1: begin
          if(_mul_12_source_start && _mul_12_stream_oready) begin
            _mul_12_source_start <= 0;
            _mul_12_source_busy <= 1;
          end 
          if(_mul_12_source_start && _mul_12_stream_oready) begin
            _mul_12_fsm <= _mul_12_fsm_2;
          end 
        end
        _mul_12_fsm_2: begin
          if(_mul_12_stream_oready) begin
            _mul_12_fsm <= _mul_12_fsm_3;
          end 
        end
        _mul_12_fsm_3: begin
          if(_mul_12_stream_oready && 1'd0) begin
            _mul_12_source_busy <= 0;
          end 
          if(_mul_12_stream_oready && 1'd0 && _mul_12_run_flag) begin
            _mul_12_source_start <= 1;
          end 
          if(_mul_12_stream_oready && 1'd0) begin
            _mul_12_fsm <= _mul_12_fsm_init;
          end 
          if(_mul_12_stream_oready && 1'd0 && _mul_12_run_flag) begin
            _mul_12_fsm <= _mul_12_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __reduce_max_13_x_source_ram_renable <= 0;
      __reduce_max_13_x_source_fifo_deq <= 0;
      __reduce_max_13_x_idle <= 1;
      __reduce_max_13_data_sink_wenable <= 0;
      __reduce_max_13_data_sink_fifo_enq <= 0;
      __reduce_max_13_valid_sink_wenable <= 0;
      __reduce_max_13_valid_sink_fifo_enq <= 0;
      ___reduce_max_13_stream_ivalid_1 <= 0;
      _reducemax_data_272 <= -33'sd2147483648;
      _reducemax_count_272 <= 0;
      _reducemax_prev_count_max_272 <= 0;
      _pulse_data_274 <= 1'sd0;
      _pulse_count_274 <= 0;
      _pulse_prev_count_max_274 <= 0;
      __variable_wdata_271 <= 0;
      __variable_wdata_269 <= 0;
      __variable_wdata_270 <= 0;
      _tmp_996 <= 0;
      _tmp_997 <= 0;
      _tmp_998 <= 0;
      _tmp_999 <= 0;
      _tmp_1000 <= 0;
      _tmp_1001 <= 0;
      _tmp_1002 <= 0;
      _tmp_1003 <= 0;
      _tmp_1004 <= 0;
      _tmp_1005 <= 0;
      _tmp_1006 <= 0;
      _tmp_1007 <= 0;
      _tmp_1008 <= 0;
      _tmp_1009 <= 0;
      _tmp_1010 <= 0;
      _tmp_1011 <= 0;
      _tmp_1012 <= 0;
      _tmp_1013 <= 0;
      _tmp_1014 <= 0;
      _tmp_1015 <= 0;
      __reduce_max_13_busy_reg <= 0;
    end else begin
      if(__reduce_max_13_stream_oready) begin
        __reduce_max_13_x_source_ram_renable <= 0;
        __reduce_max_13_x_source_fifo_deq <= 0;
      end 
      __reduce_max_13_x_idle <= __reduce_max_13_x_idle;
      if(__reduce_max_13_stream_oready) begin
        __reduce_max_13_data_sink_wenable <= 0;
        __reduce_max_13_data_sink_fifo_enq <= 0;
      end 
      if(__reduce_max_13_stream_oready) begin
        __reduce_max_13_valid_sink_wenable <= 0;
        __reduce_max_13_valid_sink_fifo_enq <= 0;
      end 
      if(__reduce_max_13_stream_oready) begin
        ___reduce_max_13_stream_ivalid_1 <= __reduce_max_13_stream_ivalid;
      end 
      if(__reduce_max_13_stream_ivalid && __reduce_max_13_stream_oready && _reducemax_reset_cond_272) begin
        _reducemax_data_272 <= -33'sd2147483648;
      end 
      if(__reduce_max_13_stream_ivalid && __reduce_max_13_stream_oready) begin
        _reducemax_count_272 <= (_reducemax_current_count_272 >= _reduce_max_13_size_data - 1)? 0 : _reducemax_current_count_272 + 1;
      end 
      if(__reduce_max_13_stream_ivalid && __reduce_max_13_stream_oready) begin
        _reducemax_prev_count_max_272 <= _reducemax_current_count_272 >= _reduce_max_13_size_data - 1;
      end 
      if(__reduce_max_13_stream_ivalid && __reduce_max_13_stream_oready) begin
        _reducemax_data_272 <= (_reducemax_current_data_272 < _reduce_max_13_x_data)? _reduce_max_13_x_data : _reducemax_current_data_272;
      end 
      if(__reduce_max_13_stream_ivalid && __reduce_max_13_stream_oready && _pulse_reset_cond_274) begin
        _pulse_data_274 <= 1'sd0;
      end 
      if(__reduce_max_13_stream_ivalid && __reduce_max_13_stream_oready) begin
        _pulse_count_274 <= (_pulse_current_count_274 >= _reduce_max_13_size_data - 1)? 0 : _pulse_current_count_274 + 1;
      end 
      if(__reduce_max_13_stream_ivalid && __reduce_max_13_stream_oready) begin
        _pulse_prev_count_max_274 <= _pulse_current_count_274 >= _reduce_max_13_size_data - 1;
      end 
      if(__reduce_max_13_stream_ivalid && __reduce_max_13_stream_oready) begin
        _pulse_data_274 <= _pulse_current_count_274 >= _reduce_max_13_size_data - 1;
      end 
      if(__stream_max_pool_serial_27_stream_ivalid_3 && _stream_max_pool_serial_27_stream_oready) begin
        __variable_wdata_271 <= __delay_data_1128__delay_1127__delay_1126__variable_883;
      end 
      if(__stream_max_pool_serial_27_stream_ivalid_3 && _stream_max_pool_serial_27_stream_oready) begin
        __variable_wdata_269 <= _cond_data_894;
      end 
      if(__stream_max_pool_serial_27_stream_ivalid_3 && _stream_max_pool_serial_27_stream_oready) begin
        __variable_wdata_270 <= __delay_data_1131__delay_1130__delay_1129__variable_880;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_996 <= __reduce_max_13_source_start;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_997 <= _tmp_996;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_998 <= _tmp_997;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_999 <= __reduce_max_13_source_start;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_1000 <= _tmp_999;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_1001 <= _tmp_1000;
      end 
      if(__reduce_max_13_stream_oready && _tmp_1001) begin
        __variable_wdata_271 <= 1;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_1002 <= __reduce_max_13_source_start;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_1003 <= _tmp_1002;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_1004 <= _tmp_1003;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_1005 <= _tmp_1004;
      end 
      if(__reduce_max_13_stream_oready && _tmp_1005) begin
        __variable_wdata_271 <= 0;
      end 
      if(__reduce_max_13_stream_oready && 1'd0) begin
        __variable_wdata_271 <= 1;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_1006 <= __reduce_max_13_source_start;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_1007 <= _tmp_1006;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_1008 <= _tmp_1007;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_1009 <= __reduce_max_13_source_stop;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_1010 <= _tmp_1009;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_1011 <= _tmp_1010;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_1012 <= __reduce_max_13_source_busy;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_1013 <= _tmp_1012;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_1014 <= _tmp_1013;
      end 
      if(__reduce_max_13_stream_oready) begin
        _tmp_1015 <= __reduce_max_13_sink_busy;
      end 
      if(!__reduce_max_13_sink_busy && _tmp_1015) begin
        __reduce_max_13_busy_reg <= 0;
      end 
      if(__reduce_max_13_source_busy) begin
        __reduce_max_13_busy_reg <= 1;
      end 
    end
  end

  localparam __reduce_max_13_fsm_1 = 1;
  localparam __reduce_max_13_fsm_2 = 2;
  localparam __reduce_max_13_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      __reduce_max_13_fsm <= __reduce_max_13_fsm_init;
      __reduce_max_13_source_start <= 0;
      __reduce_max_13_source_busy <= 0;
      __reduce_max_13_stream_ivalid <= 0;
    end else begin
      if(__stream_max_pool_serial_27_stream_ivalid_3 && _stream_max_pool_serial_27_stream_oready) begin
        __reduce_max_13_stream_ivalid <= 1'd1;
      end 
      if(_stream_max_pool_serial_27_stream_oready && _stream_max_pool_serial_27_busy) begin
        __reduce_max_13_source_busy <= _stream_max_pool_serial_27_source_busy;
      end 
      if(__reduce_max_13_stream_oready && _tmp_998) begin
        __reduce_max_13_stream_ivalid <= 1;
      end 
      if(__reduce_max_13_stream_oready && 1'd0) begin
        __reduce_max_13_stream_ivalid <= 0;
      end 
      case(__reduce_max_13_fsm)
        __reduce_max_13_fsm_init: begin
          if(__reduce_max_13_run_flag) begin
            __reduce_max_13_source_start <= 1;
          end 
          if(__reduce_max_13_run_flag) begin
            __reduce_max_13_fsm <= __reduce_max_13_fsm_1;
          end 
        end
        __reduce_max_13_fsm_1: begin
          if(__reduce_max_13_source_start && __reduce_max_13_stream_oready) begin
            __reduce_max_13_source_start <= 0;
            __reduce_max_13_source_busy <= 1;
          end 
          if(__reduce_max_13_source_start && __reduce_max_13_stream_oready) begin
            __reduce_max_13_fsm <= __reduce_max_13_fsm_2;
          end 
        end
        __reduce_max_13_fsm_2: begin
          if(__reduce_max_13_stream_oready) begin
            __reduce_max_13_fsm <= __reduce_max_13_fsm_3;
          end 
        end
        __reduce_max_13_fsm_3: begin
          if(__reduce_max_13_stream_oready && 1'd0) begin
            __reduce_max_13_source_busy <= 0;
          end 
          if(__reduce_max_13_stream_oready && 1'd0 && __reduce_max_13_run_flag) begin
            __reduce_max_13_source_start <= 1;
          end 
          if(__reduce_max_13_stream_oready && 1'd0) begin
            __reduce_max_13_fsm <= __reduce_max_13_fsm_init;
          end 
          if(__reduce_max_13_stream_oready && 1'd0 && __reduce_max_13_run_flag) begin
            __reduce_max_13_fsm <= __reduce_max_13_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_7_source_ram_renable <= 0;
      _stream_conv2d_25_source_7_source_fifo_deq <= 0;
      _stream_conv2d_25_source_7_idle <= 1;
      _stream_conv2d_25_source_9_source_ram_renable <= 0;
      _stream_conv2d_25_source_9_source_fifo_deq <= 0;
      _stream_conv2d_25_source_9_idle <= 1;
      _stream_conv2d_25_source_11_source_ram_renable <= 0;
      _stream_conv2d_25_source_11_source_fifo_deq <= 0;
      _stream_conv2d_25_source_11_idle <= 1;
      _stream_conv2d_25_source_13_source_ram_renable <= 0;
      _stream_conv2d_25_source_13_source_fifo_deq <= 0;
      _stream_conv2d_25_source_13_idle <= 1;
      _stream_conv2d_25_source_15_source_ram_renable <= 0;
      _stream_conv2d_25_source_15_source_fifo_deq <= 0;
      _stream_conv2d_25_source_15_idle <= 1;
      _stream_conv2d_25_source_20_source_ram_renable <= 0;
      _stream_conv2d_25_source_20_source_fifo_deq <= 0;
      _stream_conv2d_25_source_20_idle <= 1;
      _stream_conv2d_25_source_21_source_ram_renable <= 0;
      _stream_conv2d_25_source_21_source_fifo_deq <= 0;
      _stream_conv2d_25_source_21_idle <= 1;
      _stream_conv2d_25_source_22_source_ram_renable <= 0;
      _stream_conv2d_25_source_22_source_fifo_deq <= 0;
      _stream_conv2d_25_source_22_idle <= 1;
      _stream_conv2d_25_source_23_source_ram_renable <= 0;
      _stream_conv2d_25_source_23_source_fifo_deq <= 0;
      _stream_conv2d_25_source_23_idle <= 1;
      _stream_conv2d_25_source_24_source_ram_renable <= 0;
      _stream_conv2d_25_source_24_source_fifo_deq <= 0;
      _stream_conv2d_25_source_24_idle <= 1;
      _stream_conv2d_25_source_25_source_ram_renable <= 0;
      _stream_conv2d_25_source_25_source_fifo_deq <= 0;
      _stream_conv2d_25_source_25_idle <= 1;
      _stream_conv2d_25_source_26_source_ram_renable <= 0;
      _stream_conv2d_25_source_26_source_fifo_deq <= 0;
      _stream_conv2d_25_source_26_idle <= 1;
      _stream_conv2d_25_source_27_source_ram_renable <= 0;
      _stream_conv2d_25_source_27_source_fifo_deq <= 0;
      _stream_conv2d_25_source_27_idle <= 1;
      _stream_conv2d_25_source_28_source_ram_renable <= 0;
      _stream_conv2d_25_source_28_source_fifo_deq <= 0;
      _stream_conv2d_25_source_28_idle <= 1;
      _stream_conv2d_25_source_29_source_ram_renable <= 0;
      _stream_conv2d_25_source_29_source_fifo_deq <= 0;
      _stream_conv2d_25_source_29_idle <= 1;
      _stream_conv2d_25_source_30_source_ram_renable <= 0;
      _stream_conv2d_25_source_30_source_fifo_deq <= 0;
      _stream_conv2d_25_source_30_idle <= 1;
      _stream_conv2d_25_source_31_source_ram_renable <= 0;
      _stream_conv2d_25_source_31_source_fifo_deq <= 0;
      _stream_conv2d_25_source_31_idle <= 1;
      _stream_conv2d_25_source_32_source_ram_renable <= 0;
      _stream_conv2d_25_source_32_source_fifo_deq <= 0;
      _stream_conv2d_25_source_32_idle <= 1;
      _stream_conv2d_25_source_33_source_ram_renable <= 0;
      _stream_conv2d_25_source_33_source_fifo_deq <= 0;
      _stream_conv2d_25_source_33_idle <= 1;
      _stream_conv2d_25_source_34_source_ram_renable <= 0;
      _stream_conv2d_25_source_34_source_fifo_deq <= 0;
      _stream_conv2d_25_source_34_idle <= 1;
      _stream_conv2d_25_source_35_source_ram_renable <= 0;
      _stream_conv2d_25_source_35_source_fifo_deq <= 0;
      _stream_conv2d_25_source_35_idle <= 1;
      _stream_conv2d_25_source_36_source_ram_renable <= 0;
      _stream_conv2d_25_source_36_source_fifo_deq <= 0;
      _stream_conv2d_25_source_36_idle <= 1;
      _stream_conv2d_25_source_37_source_ram_renable <= 0;
      _stream_conv2d_25_source_37_source_fifo_deq <= 0;
      _stream_conv2d_25_source_37_idle <= 1;
      _stream_conv2d_25_sink_50_sink_wenable <= 0;
      _stream_conv2d_25_sink_50_sink_fifo_enq <= 0;
      _stream_conv2d_25_sink_51_sink_wenable <= 0;
      _stream_conv2d_25_sink_51_sink_fifo_enq <= 0;
      __stream_conv2d_25_stream_ivalid_1 <= 0;
      __stream_conv2d_25_stream_ivalid_2 <= 0;
      __stream_conv2d_25_stream_ivalid_3 <= 0;
      __stream_conv2d_25_stream_ivalid_4 <= 0;
      __stream_conv2d_25_stream_ivalid_5 <= 0;
      __stream_conv2d_25_stream_ivalid_6 <= 0;
      __stream_conv2d_25_stream_ivalid_7 <= 0;
      __stream_conv2d_25_stream_ivalid_8 <= 0;
      __stream_conv2d_25_stream_ivalid_9 <= 0;
      __stream_conv2d_25_stream_ivalid_10 <= 0;
      __stream_conv2d_25_stream_ivalid_11 <= 0;
      __stream_conv2d_25_stream_ivalid_12 <= 0;
      __stream_conv2d_25_stream_ivalid_13 <= 0;
      __stream_conv2d_25_stream_ivalid_14 <= 0;
      __stream_conv2d_25_stream_ivalid_15 <= 0;
      __stream_conv2d_25_stream_ivalid_16 <= 0;
      __stream_conv2d_25_stream_ivalid_17 <= 0;
      __stream_conv2d_25_stream_ivalid_18 <= 0;
      __stream_conv2d_25_stream_ivalid_19 <= 0;
      __stream_conv2d_25_stream_ivalid_20 <= 0;
      __stream_conv2d_25_stream_ivalid_21 <= 0;
      __stream_conv2d_25_stream_ivalid_22 <= 0;
      __stream_conv2d_25_stream_ivalid_23 <= 0;
      __stream_conv2d_25_stream_ivalid_24 <= 0;
      __stream_conv2d_25_stream_ivalid_25 <= 0;
      __stream_conv2d_25_stream_ivalid_26 <= 0;
      __stream_conv2d_25_stream_ivalid_27 <= 0;
      __stream_conv2d_25_stream_ivalid_28 <= 0;
      __stream_conv2d_25_stream_ivalid_29 <= 0;
      __stream_conv2d_25_stream_ivalid_30 <= 0;
      __stream_conv2d_25_stream_ivalid_31 <= 0;
      __stream_conv2d_25_stream_ivalid_32 <= 0;
      __stream_conv2d_25_stream_ivalid_33 <= 0;
      __stream_conv2d_25_stream_ivalid_34 <= 0;
      _eq_data_339 <= 0;
      _eq_data_343 <= 0;
      _eq_data_346 <= 0;
      _eq_data_349 <= 0;
      _eq_data_353 <= 0;
      _eq_data_356 <= 0;
      _eq_data_359 <= 0;
      _eq_data_363 <= 0;
      _eq_data_366 <= 0;
      _eq_data_369 <= 0;
      _eq_data_373 <= 0;
      _eq_data_376 <= 0;
      _eq_data_379 <= 0;
      _eq_data_383 <= 0;
      _eq_data_386 <= 0;
      _eq_data_389 <= 0;
      _eq_data_393 <= 0;
      _eq_data_396 <= 0;
      _eq_data_399 <= 0;
      _eq_data_403 <= 0;
      _eq_data_406 <= 0;
      _eq_data_409 <= 0;
      _eq_data_413 <= 0;
      _eq_data_416 <= 0;
      _eq_data_419 <= 0;
      _eq_data_423 <= 0;
      _eq_data_426 <= 0;
      _eq_data_429 <= 0;
      _eq_data_433 <= 0;
      _eq_data_436 <= 0;
      _eq_data_439 <= 0;
      _eq_data_443 <= 0;
      _eq_data_446 <= 0;
      _eq_data_449 <= 0;
      _eq_data_453 <= 0;
      _eq_data_456 <= 0;
      _eq_data_459 <= 0;
      _eq_data_463 <= 0;
      _eq_data_466 <= 0;
      _eq_data_469 <= 0;
      _eq_data_473 <= 0;
      _eq_data_476 <= 0;
      _eq_data_479 <= 0;
      _eq_data_483 <= 0;
      _eq_data_486 <= 0;
      _eq_data_489 <= 0;
      _eq_data_493 <= 0;
      _eq_data_496 <= 0;
      _eq_data_499 <= 0;
      _eq_data_503 <= 0;
      _eq_data_506 <= 0;
      _eq_data_509 <= 0;
      _eq_data_513 <= 0;
      _eq_data_516 <= 0;
      _plus_data_671 <= 0;
      _plus_data_690 <= 0;
      _plus_data_709 <= 0;
      _plus_data_728 <= 0;
      _plus_data_747 <= 0;
      _plus_data_766 <= 0;
      _plus_data_785 <= 0;
      _plus_data_804 <= 0;
      _plus_data_823 <= 0;
      _plus_data_839 <= 0;
      _plus_data_858 <= 0;
      __delay_data_946__variable_332 <= 0;
      __delay_data_947__variable_331 <= 0;
      __delay_data_948__variable_330 <= 0;
      __delay_data_949__variable_335 <= 0;
      __delay_data_950__variable_334 <= 0;
      __delay_data_951__variable_333 <= 0;
      __delay_data_952__variable_338 <= 0;
      __delay_data_953__variable_337 <= 0;
      __delay_data_954__variable_336 <= 0;
      __delay_data_955_pointer_618 <= 0;
      __delay_data_956_reinterpretcast_609 <= 0;
      __delay_data_957_pointer_620 <= 0;
      __delay_data_958_reinterpretcast_610 <= 0;
      __delay_data_959_pointer_622 <= 0;
      __delay_data_960_reinterpretcast_611 <= 0;
      __delay_data_961_pointer_624 <= 0;
      __delay_data_962_reinterpretcast_612 <= 0;
      __delay_data_963_pointer_626 <= 0;
      __delay_data_964_reinterpretcast_613 <= 0;
      __delay_data_965_pointer_628 <= 0;
      __delay_data_966_reinterpretcast_614 <= 0;
      __delay_data_967_pointer_630 <= 0;
      __delay_data_968_reinterpretcast_615 <= 0;
      __delay_data_969_pointer_632 <= 0;
      __delay_data_970_reinterpretcast_616 <= 0;
      __delay_data_971_pointer_634 <= 0;
      __delay_data_972_reinterpretcast_617 <= 0;
      __delay_data_973__variable_281 <= 0;
      __delay_data_998__variable_276 <= 0;
      __delay_data_1011_cond_297 <= 0;
      __delay_data_1030_cond_304 <= 0;
      __delay_data_1069_eq_873 <= 0;
      __delay_data_974__delay_973__variable_281 <= 0;
      __delay_data_986_plus_839 <= 0;
      __delay_data_999__delay_998__variable_276 <= 0;
      __delay_data_1012__delay_1011_cond_297 <= 0;
      __delay_data_1031__delay_1030_cond_304 <= 0;
      __delay_data_1050_plus_858 <= 0;
      __delay_data_1070__delay_1069_eq_873 <= 0;
      __delay_data_975__delay_974__delay_973__variable_281 <= 0;
      __delay_data_987__delay_986_plus_839 <= 0;
      __delay_data_1000__delay_999__delay_998__variable_276 <= 0;
      __delay_data_1013__delay_1012__delay_1011_cond_297 <= 0;
      __delay_data_1032__delay_1031__delay_1030_cond_304 <= 0;
      __delay_data_1051__delay_1050_plus_858 <= 0;
      __delay_data_1071__delay_1070__delay_1069_eq_873 <= 0;
      __delay_data_976__delay_975__delay_974____variable_281 <= 0;
      __delay_data_988__delay_987__delay_986_plus_839 <= 0;
      __delay_data_1001__delay_1000__delay_999____variable_276 <= 0;
      __delay_data_1014__delay_1013__delay_1012__delay_1011_cond_297 <= 0;
      __delay_data_1033__delay_1032__delay_1031__delay_1030_cond_304 <= 0;
      __delay_data_1052__delay_1051__delay_1050_plus_858 <= 0;
      __delay_data_1072__delay_1071__delay_1070__delay_1069_eq_873 <= 0;
      __delay_data_977__delay_976__delay_975____variable_281 <= 0;
      __delay_data_989__delay_988__delay_987__delay_986_plus_839 <= 0;
      __delay_data_1002__delay_1001__delay_1000____variable_276 <= 0;
      __delay_data_1015__delay_1014__delay_1013__delay_1012___cond_297 <= 0;
      __delay_data_1034__delay_1033__delay_1032__delay_1031___cond_304 <= 0;
      __delay_data_1053__delay_1052__delay_1051__delay_1050_plus_858 <= 0;
      __delay_data_1073__delay_1072__delay_1071__delay_1070___eq_873 <= 0;
      __delay_data_978__delay_977__delay_976____variable_281 <= 0;
      __delay_data_990__delay_989__delay_988__delay_987___plus_839 <= 0;
      __delay_data_1003__delay_1002__delay_1001____variable_276 <= 0;
      __delay_data_1016__delay_1015__delay_1014__delay_1013___cond_297 <= 0;
      __delay_data_1035__delay_1034__delay_1033__delay_1032___cond_304 <= 0;
      __delay_data_1054__delay_1053__delay_1052__delay_1051___plus_858 <= 0;
      __delay_data_1074__delay_1073__delay_1072__delay_1071___eq_873 <= 0;
      __delay_data_979__delay_978__delay_977____variable_281 <= 0;
      __delay_data_991__delay_990__delay_989__delay_988___plus_839 <= 0;
      __delay_data_1004__delay_1003__delay_1002____variable_276 <= 0;
      __delay_data_1017__delay_1016__delay_1015__delay_1014___cond_297 <= 0;
      __delay_data_1036__delay_1035__delay_1034__delay_1033___cond_304 <= 0;
      __delay_data_1055__delay_1054__delay_1053__delay_1052___plus_858 <= 0;
      __delay_data_1075__delay_1074__delay_1073__delay_1072___eq_873 <= 0;
      __delay_data_980__delay_979__delay_978____variable_281 <= 0;
      __delay_data_992__delay_991__delay_990__delay_989___plus_839 <= 0;
      __delay_data_1005__delay_1004__delay_1003____variable_276 <= 0;
      __delay_data_1018__delay_1017__delay_1016__delay_1015___cond_297 <= 0;
      __delay_data_1037__delay_1036__delay_1035__delay_1034___cond_304 <= 0;
      __delay_data_1056__delay_1055__delay_1054__delay_1053___plus_858 <= 0;
      __delay_data_1076__delay_1075__delay_1074__delay_1073___eq_873 <= 0;
      __delay_data_981__delay_980__delay_979____variable_281 <= 0;
      __delay_data_993__delay_992__delay_991__delay_990___plus_839 <= 0;
      __delay_data_1006__delay_1005__delay_1004____variable_276 <= 0;
      __delay_data_1019__delay_1018__delay_1017__delay_1016___cond_297 <= 0;
      __delay_data_1038__delay_1037__delay_1036__delay_1035___cond_304 <= 0;
      __delay_data_1057__delay_1056__delay_1055__delay_1054___plus_858 <= 0;
      __delay_data_1077__delay_1076__delay_1075__delay_1074___eq_873 <= 0;
      __delay_data_982__delay_981__delay_980____variable_281 <= 0;
      __delay_data_994__delay_993__delay_992__delay_991___plus_839 <= 0;
      __delay_data_1007__delay_1006__delay_1005____variable_276 <= 0;
      __delay_data_1020__delay_1019__delay_1018__delay_1017___cond_297 <= 0;
      __delay_data_1039__delay_1038__delay_1037__delay_1036___cond_304 <= 0;
      __delay_data_1058__delay_1057__delay_1056__delay_1055___plus_858 <= 0;
      __delay_data_1078__delay_1077__delay_1076__delay_1075___eq_873 <= 0;
      __delay_data_983__delay_982__delay_981____variable_281 <= 0;
      __delay_data_995__delay_994__delay_993__delay_992___plus_839 <= 0;
      __delay_data_1008__delay_1007__delay_1006____variable_276 <= 0;
      __delay_data_1021__delay_1020__delay_1019__delay_1018___cond_297 <= 0;
      __delay_data_1040__delay_1039__delay_1038__delay_1037___cond_304 <= 0;
      __delay_data_1059__delay_1058__delay_1057__delay_1056___plus_858 <= 0;
      __delay_data_1079__delay_1078__delay_1077__delay_1076___eq_873 <= 0;
      __delay_data_984__delay_983__delay_982____variable_281 <= 0;
      __delay_data_996__delay_995__delay_994__delay_993___plus_839 <= 0;
      __delay_data_1009__delay_1008__delay_1007____variable_276 <= 0;
      __delay_data_1022__delay_1021__delay_1020__delay_1019___cond_297 <= 0;
      __delay_data_1041__delay_1040__delay_1039__delay_1038___cond_304 <= 0;
      __delay_data_1060__delay_1059__delay_1058__delay_1057___plus_858 <= 0;
      __delay_data_1080__delay_1079__delay_1078__delay_1077___eq_873 <= 0;
      __delay_data_985__delay_984__delay_983____variable_281 <= 0;
      __delay_data_997__delay_996__delay_995__delay_994___plus_839 <= 0;
      __delay_data_1010__delay_1009__delay_1008____variable_276 <= 0;
      __delay_data_1023__delay_1022__delay_1021__delay_1020___cond_297 <= 0;
      __delay_data_1042__delay_1041__delay_1040__delay_1039___cond_304 <= 0;
      __delay_data_1061__delay_1060__delay_1059__delay_1058___plus_858 <= 0;
      __delay_data_1081__delay_1080__delay_1079__delay_1078___eq_873 <= 0;
      __delay_data_1024__delay_1023__delay_1022__delay_1021___cond_297 <= 0;
      __delay_data_1043__delay_1042__delay_1041__delay_1040___cond_304 <= 0;
      __delay_data_1062__delay_1061__delay_1060__delay_1059___plus_858 <= 0;
      __delay_data_1082__delay_1081__delay_1080__delay_1079___eq_873 <= 0;
      __delay_data_1025__delay_1024__delay_1023__delay_1022___cond_297 <= 0;
      __delay_data_1044__delay_1043__delay_1042__delay_1041___cond_304 <= 0;
      __delay_data_1063__delay_1062__delay_1061__delay_1060___plus_858 <= 0;
      __delay_data_1083__delay_1082__delay_1081__delay_1080___eq_873 <= 0;
      __delay_data_1026__delay_1025__delay_1024__delay_1023___cond_297 <= 0;
      __delay_data_1045__delay_1044__delay_1043__delay_1042___cond_304 <= 0;
      __delay_data_1064__delay_1063__delay_1062__delay_1061___plus_858 <= 0;
      __delay_data_1084__delay_1083__delay_1082__delay_1081___eq_873 <= 0;
      __delay_data_1027__delay_1026__delay_1025__delay_1024___cond_297 <= 0;
      __delay_data_1046__delay_1045__delay_1044__delay_1043___cond_304 <= 0;
      __delay_data_1065__delay_1064__delay_1063__delay_1062___plus_858 <= 0;
      __delay_data_1085__delay_1084__delay_1083__delay_1082___eq_873 <= 0;
      __delay_data_1028__delay_1027__delay_1026__delay_1025___cond_297 <= 0;
      __delay_data_1047__delay_1046__delay_1045__delay_1044___cond_304 <= 0;
      __delay_data_1066__delay_1065__delay_1064__delay_1063___plus_858 <= 0;
      __delay_data_1086__delay_1085__delay_1084__delay_1083___eq_873 <= 0;
      __delay_data_1029__delay_1028__delay_1027__delay_1026___cond_297 <= 0;
      __delay_data_1048__delay_1047__delay_1046__delay_1045___cond_304 <= 0;
      __delay_data_1067__delay_1066__delay_1065__delay_1064___plus_858 <= 0;
      __delay_data_1087__delay_1086__delay_1085__delay_1084___eq_873 <= 0;
      _plus_data_842 <= 0;
      __delay_data_1049__delay_1048__delay_1047__delay_1046___cond_304 <= 0;
      __delay_data_1068__delay_1067__delay_1066__delay_1065___plus_858 <= 0;
      __delay_data_1088__delay_1087__delay_1086__delay_1085___eq_873 <= 0;
      __delay_data_1108__substreamoutput_841 <= 0;
      __delay_data_1089__delay_1088__delay_1087__delay_1086___eq_873 <= 0;
      __delay_data_1109__delay_1108__substreamoutput_841 <= 0;
      __delay_data_1090__delay_1089__delay_1088__delay_1087___eq_873 <= 0;
      __delay_data_1110__delay_1109__delay_1108__substreamoutput_841 <= 0;
      __delay_data_1091__delay_1090__delay_1089__delay_1088___eq_873 <= 0;
      __delay_data_1111__delay_1110__delay_1109____substreamoutput_841 <= 0;
      __delay_data_1092__delay_1091__delay_1090__delay_1089___eq_873 <= 0;
      __delay_data_1112__delay_1111__delay_1110____substreamoutput_841 <= 0;
      __delay_data_1093__delay_1092__delay_1091__delay_1090___eq_873 <= 0;
      __delay_data_1113__delay_1112__delay_1111____substreamoutput_841 <= 0;
      __delay_data_1094__delay_1093__delay_1092__delay_1091___eq_873 <= 0;
      __delay_data_1114__delay_1113__delay_1112____substreamoutput_841 <= 0;
      __delay_data_1095__delay_1094__delay_1093__delay_1092___eq_873 <= 0;
      __delay_data_1115__delay_1114__delay_1113____substreamoutput_841 <= 0;
      __delay_data_1096__delay_1095__delay_1094__delay_1093___eq_873 <= 0;
      __delay_data_1116__delay_1115__delay_1114____substreamoutput_841 <= 0;
      __delay_data_1097__delay_1096__delay_1095__delay_1094___eq_873 <= 0;
      __delay_data_1117__delay_1116__delay_1115____substreamoutput_841 <= 0;
      _times_mul_odata_reg_860 <= 0;
      _greaterthan_data_877 <= 0;
      __delay_data_1098__delay_1097__delay_1096__delay_1095___eq_873 <= 0;
      __delay_data_1104__substreamoutput_859 <= 0;
      __delay_data_1118__delay_1117__delay_1116____substreamoutput_841 <= 0;
      __delay_data_1099__delay_1098__delay_1097__delay_1096___eq_873 <= 0;
      __delay_data_1101_greaterthan_877 <= 0;
      __delay_data_1105__delay_1104__substreamoutput_859 <= 0;
      __delay_data_1119__delay_1118__delay_1117____substreamoutput_841 <= 0;
      __delay_data_1100__delay_1099__delay_1098__delay_1097___eq_873 <= 0;
      __delay_data_1102__delay_1101_greaterthan_877 <= 0;
      __delay_data_1106__delay_1105__delay_1104__substreamoutput_859 <= 0;
      __delay_data_1120__delay_1119__delay_1118____substreamoutput_841 <= 0;
      _cond_data_875 <= 0;
      __delay_data_1103__delay_1102__delay_1101_greaterthan_877 <= 0;
      __delay_data_1107__delay_1106__delay_1105____substreamoutput_859 <= 0;
      __delay_data_1121__delay_1120__delay_1119____substreamoutput_841 <= 0;
      _cond_data_878 <= 0;
      __delay_data_1122__delay_1121__delay_1120____substreamoutput_841 <= 0;
      _stream_conv2d_25_parameter_0_next_parameter_data <= 0;
      __variable_wdata_276 <= 0;
      _stream_conv2d_25_parameter_1_next_parameter_data <= 0;
      __variable_wdata_277 <= 0;
      _stream_conv2d_25_parameter_2_next_parameter_data <= 0;
      __variable_wdata_278 <= 0;
      _stream_conv2d_25_parameter_3_next_parameter_data <= 0;
      __variable_wdata_279 <= 0;
      _stream_conv2d_25_parameter_4_next_parameter_data <= 0;
      __variable_wdata_280 <= 0;
      _stream_conv2d_25_parameter_6_next_parameter_data <= 0;
      __variable_wdata_291 <= 0;
      _stream_conv2d_25_source_7_source_mode <= 5'b0;
      _stream_conv2d_25_source_7_source_offset <= 0;
      _source_stream_conv2d_25_source_7_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_7_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_7_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_7_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_7_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_7_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_7_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_7_pat_stride_3 <= 0;
      _stream_conv2d_25_source_7_source_sel <= 0;
      _stream_conv2d_25_source_7_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_7_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_7_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_7_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_7_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_7_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_7_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_7_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_7_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_7_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_7_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_7_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_7_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_7_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_7_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_7_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_7_pat_stride_buf_3 <= 0;
      __variable_wdata_292 <= 0;
      _stream_conv2d_25_source_7_source_ram_raddr <= 0;
      _stream_conv2d_25_parameter_8_next_parameter_data <= 0;
      __variable_wdata_298 <= 0;
      _stream_conv2d_25_source_9_source_mode <= 5'b0;
      _stream_conv2d_25_source_9_source_offset <= 0;
      _source_stream_conv2d_25_source_9_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_9_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_9_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_9_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_9_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_9_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_9_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_9_pat_stride_3 <= 0;
      _stream_conv2d_25_source_9_source_sel <= 0;
      _stream_conv2d_25_source_9_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_9_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_9_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_9_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_9_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_9_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_9_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_9_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_9_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_9_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_9_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_9_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_9_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_9_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_9_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_9_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_9_pat_stride_buf_3 <= 0;
      __variable_wdata_299 <= 0;
      _stream_conv2d_25_source_9_source_ram_raddr <= 0;
      _stream_conv2d_25_parameter_10_next_parameter_data <= 0;
      __variable_wdata_305 <= 0;
      _stream_conv2d_25_source_11_source_mode <= 5'b0;
      _stream_conv2d_25_source_11_source_empty_data <= 0;
      __variable_wdata_306 <= 0;
      _stream_conv2d_25_parameter_12_next_parameter_data <= 0;
      __variable_wdata_312 <= 0;
      _stream_conv2d_25_source_13_source_mode <= 5'b0;
      _stream_conv2d_25_source_13_source_empty_data <= 0;
      __variable_wdata_313 <= 0;
      _stream_conv2d_25_parameter_14_next_parameter_data <= 0;
      __variable_wdata_319 <= 0;
      _stream_conv2d_25_source_15_source_mode <= 5'b0;
      _stream_conv2d_25_source_15_source_empty_data <= 0;
      __variable_wdata_320 <= 0;
      _stream_conv2d_25_parameter_16_next_parameter_data <= 0;
      __variable_wdata_326 <= 0;
      _stream_conv2d_25_parameter_17_next_parameter_data <= 0;
      __variable_wdata_327 <= 0;
      _stream_conv2d_25_parameter_18_next_parameter_data <= 0;
      __variable_wdata_328 <= 0;
      _stream_conv2d_25_parameter_19_next_parameter_data <= 0;
      __variable_wdata_329 <= 0;
      _stream_conv2d_25_source_20_source_mode <= 5'b0;
      _stream_conv2d_25_source_20_source_offset <= 0;
      _source_stream_conv2d_25_source_20_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_20_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_20_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_20_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_20_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_20_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_20_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_20_pat_stride_3 <= 0;
      _stream_conv2d_25_source_20_source_sel <= 0;
      _stream_conv2d_25_source_20_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_20_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_20_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_20_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_20_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_20_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_20_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_20_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_20_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_20_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_20_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_20_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_20_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_20_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_20_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_20_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_20_pat_stride_buf_3 <= 0;
      __variable_wdata_330 <= 0;
      _stream_conv2d_25_source_20_source_ram_raddr <= 0;
      _stream_conv2d_25_source_21_source_mode <= 5'b0;
      _stream_conv2d_25_source_21_source_offset <= 0;
      _source_stream_conv2d_25_source_21_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_21_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_21_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_21_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_21_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_21_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_21_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_21_pat_stride_3 <= 0;
      _stream_conv2d_25_source_21_source_sel <= 0;
      _stream_conv2d_25_source_21_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_21_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_21_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_21_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_21_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_21_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_21_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_21_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_21_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_21_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_21_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_21_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_21_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_21_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_21_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_21_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_21_pat_stride_buf_3 <= 0;
      __variable_wdata_331 <= 0;
      _stream_conv2d_25_source_21_source_ram_raddr <= 0;
      _stream_conv2d_25_source_22_source_mode <= 5'b0;
      _stream_conv2d_25_source_22_source_offset <= 0;
      _source_stream_conv2d_25_source_22_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_22_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_22_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_22_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_22_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_22_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_22_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_22_pat_stride_3 <= 0;
      _stream_conv2d_25_source_22_source_sel <= 0;
      _stream_conv2d_25_source_22_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_22_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_22_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_22_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_22_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_22_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_22_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_22_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_22_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_22_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_22_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_22_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_22_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_22_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_22_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_22_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_22_pat_stride_buf_3 <= 0;
      __variable_wdata_332 <= 0;
      _stream_conv2d_25_source_22_source_ram_raddr <= 0;
      _stream_conv2d_25_source_23_source_mode <= 5'b0;
      _stream_conv2d_25_source_23_source_offset <= 0;
      _source_stream_conv2d_25_source_23_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_23_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_23_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_23_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_23_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_23_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_23_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_23_pat_stride_3 <= 0;
      _stream_conv2d_25_source_23_source_sel <= 0;
      _stream_conv2d_25_source_23_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_23_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_23_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_23_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_23_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_23_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_23_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_23_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_23_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_23_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_23_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_23_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_23_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_23_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_23_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_23_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_23_pat_stride_buf_3 <= 0;
      __variable_wdata_333 <= 0;
      _stream_conv2d_25_source_23_source_ram_raddr <= 0;
      _stream_conv2d_25_source_24_source_mode <= 5'b0;
      _stream_conv2d_25_source_24_source_offset <= 0;
      _source_stream_conv2d_25_source_24_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_24_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_24_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_24_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_24_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_24_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_24_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_24_pat_stride_3 <= 0;
      _stream_conv2d_25_source_24_source_sel <= 0;
      _stream_conv2d_25_source_24_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_24_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_24_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_24_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_24_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_24_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_24_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_24_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_24_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_24_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_24_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_24_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_24_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_24_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_24_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_24_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_24_pat_stride_buf_3 <= 0;
      __variable_wdata_334 <= 0;
      _stream_conv2d_25_source_24_source_ram_raddr <= 0;
      _stream_conv2d_25_source_25_source_mode <= 5'b0;
      _stream_conv2d_25_source_25_source_offset <= 0;
      _source_stream_conv2d_25_source_25_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_25_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_25_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_25_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_25_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_25_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_25_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_25_pat_stride_3 <= 0;
      _stream_conv2d_25_source_25_source_sel <= 0;
      _stream_conv2d_25_source_25_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_25_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_25_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_25_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_25_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_25_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_25_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_25_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_25_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_25_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_25_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_25_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_25_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_25_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_25_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_25_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_25_pat_stride_buf_3 <= 0;
      __variable_wdata_335 <= 0;
      _stream_conv2d_25_source_25_source_ram_raddr <= 0;
      _stream_conv2d_25_source_26_source_mode <= 5'b0;
      _stream_conv2d_25_source_26_source_offset <= 0;
      _source_stream_conv2d_25_source_26_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_26_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_26_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_26_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_26_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_26_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_26_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_26_pat_stride_3 <= 0;
      _stream_conv2d_25_source_26_source_sel <= 0;
      _stream_conv2d_25_source_26_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_26_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_26_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_26_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_26_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_26_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_26_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_26_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_26_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_26_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_26_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_26_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_26_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_26_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_26_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_26_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_26_pat_stride_buf_3 <= 0;
      __variable_wdata_336 <= 0;
      _stream_conv2d_25_source_26_source_ram_raddr <= 0;
      _stream_conv2d_25_source_27_source_mode <= 5'b0;
      _stream_conv2d_25_source_27_source_offset <= 0;
      _source_stream_conv2d_25_source_27_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_27_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_27_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_27_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_27_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_27_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_27_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_27_pat_stride_3 <= 0;
      _stream_conv2d_25_source_27_source_sel <= 0;
      _stream_conv2d_25_source_27_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_27_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_27_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_27_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_27_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_27_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_27_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_27_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_27_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_27_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_27_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_27_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_27_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_27_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_27_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_27_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_27_pat_stride_buf_3 <= 0;
      __variable_wdata_337 <= 0;
      _stream_conv2d_25_source_27_source_ram_raddr <= 0;
      _stream_conv2d_25_source_28_source_mode <= 5'b0;
      _stream_conv2d_25_source_28_source_offset <= 0;
      _source_stream_conv2d_25_source_28_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_28_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_28_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_28_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_28_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_28_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_28_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_28_pat_stride_3 <= 0;
      _stream_conv2d_25_source_28_source_sel <= 0;
      _stream_conv2d_25_source_28_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_28_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_28_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_28_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_28_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_28_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_28_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_28_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_28_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_28_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_28_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_28_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_28_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_28_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_28_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_28_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_28_pat_stride_buf_3 <= 0;
      __variable_wdata_338 <= 0;
      _stream_conv2d_25_source_28_source_ram_raddr <= 0;
      _stream_conv2d_25_source_29_source_mode <= 5'b0;
      _stream_conv2d_25_source_29_source_offset <= 0;
      _source_stream_conv2d_25_source_29_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_29_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_29_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_29_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_29_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_29_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_29_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_29_pat_stride_3 <= 0;
      _stream_conv2d_25_source_29_source_sel <= 0;
      _stream_conv2d_25_source_29_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_29_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_29_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_29_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_29_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_29_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_29_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_29_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_29_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_29_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_29_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_29_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_29_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_29_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_29_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_29_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_29_pat_stride_buf_3 <= 0;
      __variable_wdata_564 <= 0;
      _stream_conv2d_25_source_29_source_ram_raddr <= 0;
      _stream_conv2d_25_source_30_source_mode <= 5'b0;
      _stream_conv2d_25_source_30_source_offset <= 0;
      _source_stream_conv2d_25_source_30_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_30_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_30_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_30_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_30_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_30_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_30_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_30_pat_stride_3 <= 0;
      _stream_conv2d_25_source_30_source_sel <= 0;
      _stream_conv2d_25_source_30_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_30_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_30_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_30_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_30_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_30_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_30_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_30_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_30_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_30_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_30_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_30_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_30_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_30_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_30_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_30_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_30_pat_stride_buf_3 <= 0;
      __variable_wdata_565 <= 0;
      _stream_conv2d_25_source_30_source_ram_raddr <= 0;
      _stream_conv2d_25_source_31_source_mode <= 5'b0;
      _stream_conv2d_25_source_31_source_offset <= 0;
      _source_stream_conv2d_25_source_31_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_31_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_31_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_31_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_31_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_31_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_31_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_31_pat_stride_3 <= 0;
      _stream_conv2d_25_source_31_source_sel <= 0;
      _stream_conv2d_25_source_31_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_31_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_31_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_31_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_31_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_31_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_31_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_31_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_31_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_31_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_31_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_31_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_31_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_31_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_31_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_31_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_31_pat_stride_buf_3 <= 0;
      __variable_wdata_566 <= 0;
      _stream_conv2d_25_source_31_source_ram_raddr <= 0;
      _stream_conv2d_25_source_32_source_mode <= 5'b0;
      _stream_conv2d_25_source_32_source_offset <= 0;
      _source_stream_conv2d_25_source_32_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_32_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_32_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_32_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_32_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_32_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_32_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_32_pat_stride_3 <= 0;
      _stream_conv2d_25_source_32_source_sel <= 0;
      _stream_conv2d_25_source_32_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_32_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_32_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_32_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_32_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_32_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_32_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_32_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_32_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_32_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_32_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_32_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_32_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_32_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_32_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_32_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_32_pat_stride_buf_3 <= 0;
      __variable_wdata_567 <= 0;
      _stream_conv2d_25_source_32_source_ram_raddr <= 0;
      _stream_conv2d_25_source_33_source_mode <= 5'b0;
      _stream_conv2d_25_source_33_source_offset <= 0;
      _source_stream_conv2d_25_source_33_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_33_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_33_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_33_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_33_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_33_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_33_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_33_pat_stride_3 <= 0;
      _stream_conv2d_25_source_33_source_sel <= 0;
      _stream_conv2d_25_source_33_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_33_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_33_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_33_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_33_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_33_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_33_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_33_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_33_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_33_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_33_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_33_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_33_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_33_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_33_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_33_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_33_pat_stride_buf_3 <= 0;
      __variable_wdata_568 <= 0;
      _stream_conv2d_25_source_33_source_ram_raddr <= 0;
      _stream_conv2d_25_source_34_source_mode <= 5'b0;
      _stream_conv2d_25_source_34_source_offset <= 0;
      _source_stream_conv2d_25_source_34_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_34_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_34_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_34_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_34_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_34_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_34_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_34_pat_stride_3 <= 0;
      _stream_conv2d_25_source_34_source_sel <= 0;
      _stream_conv2d_25_source_34_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_34_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_34_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_34_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_34_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_34_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_34_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_34_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_34_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_34_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_34_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_34_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_34_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_34_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_34_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_34_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_34_pat_stride_buf_3 <= 0;
      __variable_wdata_569 <= 0;
      _stream_conv2d_25_source_34_source_ram_raddr <= 0;
      _stream_conv2d_25_source_35_source_mode <= 5'b0;
      _stream_conv2d_25_source_35_source_offset <= 0;
      _source_stream_conv2d_25_source_35_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_35_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_35_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_35_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_35_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_35_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_35_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_35_pat_stride_3 <= 0;
      _stream_conv2d_25_source_35_source_sel <= 0;
      _stream_conv2d_25_source_35_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_35_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_35_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_35_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_35_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_35_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_35_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_35_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_35_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_35_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_35_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_35_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_35_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_35_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_35_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_35_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_35_pat_stride_buf_3 <= 0;
      __variable_wdata_570 <= 0;
      _stream_conv2d_25_source_35_source_ram_raddr <= 0;
      _stream_conv2d_25_source_36_source_mode <= 5'b0;
      _stream_conv2d_25_source_36_source_offset <= 0;
      _source_stream_conv2d_25_source_36_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_36_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_36_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_36_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_36_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_36_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_36_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_36_pat_stride_3 <= 0;
      _stream_conv2d_25_source_36_source_sel <= 0;
      _stream_conv2d_25_source_36_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_36_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_36_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_36_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_36_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_36_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_36_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_36_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_36_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_36_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_36_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_36_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_36_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_36_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_36_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_36_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_36_pat_stride_buf_3 <= 0;
      __variable_wdata_571 <= 0;
      _stream_conv2d_25_source_36_source_ram_raddr <= 0;
      _stream_conv2d_25_source_37_source_mode <= 5'b0;
      _stream_conv2d_25_source_37_source_offset <= 0;
      _source_stream_conv2d_25_source_37_pat_size_0 <= 0;
      _source_stream_conv2d_25_source_37_pat_stride_0 <= 0;
      _source_stream_conv2d_25_source_37_pat_size_1 <= 0;
      _source_stream_conv2d_25_source_37_pat_stride_1 <= 0;
      _source_stream_conv2d_25_source_37_pat_size_2 <= 0;
      _source_stream_conv2d_25_source_37_pat_stride_2 <= 0;
      _source_stream_conv2d_25_source_37_pat_size_3 <= 0;
      _source_stream_conv2d_25_source_37_pat_stride_3 <= 0;
      _stream_conv2d_25_source_37_source_sel <= 0;
      _stream_conv2d_25_source_37_source_offset_buf <= 0;
      _source_stream_conv2d_25_source_37_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_25_source_37_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_25_source_37_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_25_source_37_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_25_source_37_pat_count_0 <= 0;
      _source_stream_conv2d_25_source_37_pat_count_1 <= 0;
      _source_stream_conv2d_25_source_37_pat_count_2 <= 0;
      _source_stream_conv2d_25_source_37_pat_count_3 <= 0;
      _source_stream_conv2d_25_source_37_pat_size_buf_0 <= 0;
      _source_stream_conv2d_25_source_37_pat_size_buf_1 <= 0;
      _source_stream_conv2d_25_source_37_pat_size_buf_2 <= 0;
      _source_stream_conv2d_25_source_37_pat_size_buf_3 <= 0;
      _source_stream_conv2d_25_source_37_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_25_source_37_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_25_source_37_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_25_source_37_pat_stride_buf_3 <= 0;
      __variable_wdata_572 <= 0;
      _stream_conv2d_25_source_37_source_ram_raddr <= 0;
      _tmp_296 <= 0;
      _tmp_297 <= 0;
      _tmp_298 <= 0;
      _tmp_299 <= 0;
      _tmp_300 <= 0;
      _tmp_301 <= 0;
      _tmp_302 <= 0;
      _tmp_303 <= 0;
      _tmp_304 <= 0;
      _tmp_305 <= 0;
      _tmp_306 <= 0;
      _tmp_307 <= 0;
      _tmp_308 <= 0;
      _tmp_309 <= 0;
      _tmp_310 <= 0;
      _tmp_311 <= 0;
      _tmp_312 <= 0;
      _tmp_313 <= 0;
      _tmp_314 <= 0;
      _tmp_315 <= 0;
      _tmp_316 <= 0;
      _tmp_317 <= 0;
      _tmp_318 <= 0;
      _tmp_319 <= 0;
      _tmp_320 <= 0;
      _tmp_321 <= 0;
      _tmp_322 <= 0;
      _tmp_323 <= 0;
      _tmp_324 <= 0;
      _tmp_325 <= 0;
      _tmp_326 <= 0;
      _tmp_327 <= 0;
      _tmp_328 <= 0;
      _tmp_329 <= 0;
      _tmp_330 <= 0;
      _tmp_331 <= 0;
      _tmp_334 <= 0;
      _tmp_335 <= 0;
      _tmp_336 <= 0;
      _tmp_337 <= 0;
      _tmp_338 <= 0;
      _tmp_339 <= 0;
      _tmp_340 <= 0;
      _tmp_341 <= 0;
      _tmp_342 <= 0;
      _tmp_343 <= 0;
      _tmp_344 <= 0;
      _tmp_345 <= 0;
      _tmp_346 <= 0;
      _tmp_347 <= 0;
      _tmp_348 <= 0;
      _tmp_349 <= 0;
      _tmp_350 <= 0;
      _tmp_351 <= 0;
      _tmp_352 <= 0;
      _tmp_353 <= 0;
      _tmp_354 <= 0;
      _tmp_355 <= 0;
      _tmp_356 <= 0;
      _tmp_357 <= 0;
      _tmp_358 <= 0;
      _tmp_359 <= 0;
      _tmp_360 <= 0;
      _tmp_361 <= 0;
      _tmp_362 <= 0;
      _tmp_363 <= 0;
      _tmp_364 <= 0;
      _tmp_365 <= 0;
      _tmp_366 <= 0;
      _tmp_367 <= 0;
      _tmp_368 <= 0;
      _tmp_369 <= 0;
      _tmp_370 <= 0;
      _tmp_371 <= 0;
      _tmp_372 <= 0;
      _tmp_373 <= 0;
      _tmp_374 <= 0;
      _tmp_375 <= 0;
      _tmp_376 <= 0;
      _tmp_377 <= 0;
      _tmp_378 <= 0;
      _tmp_379 <= 0;
      _tmp_380 <= 0;
      _tmp_381 <= 0;
      _tmp_382 <= 0;
      _tmp_383 <= 0;
      _tmp_384 <= 0;
      _tmp_385 <= 0;
      _tmp_386 <= 0;
      _tmp_387 <= 0;
      _tmp_388 <= 0;
      _tmp_389 <= 0;
      _tmp_390 <= 0;
      _tmp_391 <= 0;
      _tmp_392 <= 0;
      _tmp_393 <= 0;
      _tmp_394 <= 0;
      _tmp_395 <= 0;
      _tmp_396 <= 0;
      _tmp_397 <= 0;
      _tmp_398 <= 0;
      _tmp_399 <= 0;
      _tmp_400 <= 0;
      _tmp_401 <= 0;
      _tmp_402 <= 0;
      _tmp_403 <= 0;
      _tmp_404 <= 0;
      _tmp_405 <= 0;
      _stream_conv2d_25_sink_50_sink_mode <= 5'b0;
      _stream_conv2d_25_sink_50_sink_offset <= 0;
      _stream_conv2d_25_sink_50_sink_size <= 0;
      _stream_conv2d_25_sink_50_sink_stride <= 0;
      _stream_conv2d_25_sink_50_sink_sel <= 0;
      _stream_conv2d_25_sink_50_sink_offset_buf <= 0;
      _stream_conv2d_25_sink_50_sink_size_buf <= 0;
      _stream_conv2d_25_sink_50_sink_stride_buf <= 0;
      _stream_conv2d_25_sink_50_sink_waddr <= 0;
      _stream_conv2d_25_sink_50_sink_count <= 0;
      _stream_conv2d_25_sink_50_sink_wdata <= 0;
      _tmp_795 <= 0;
      _tmp_796 <= 0;
      _tmp_797 <= 0;
      _tmp_798 <= 0;
      _tmp_799 <= 0;
      _tmp_800 <= 0;
      __variable_wdata_281 <= 0;
      _tmp_801 <= 0;
      _tmp_802 <= 0;
      _tmp_803 <= 0;
      _tmp_804 <= 0;
      _tmp_807 <= 0;
      _tmp_810 <= 0;
      _tmp_811 <= 0;
      _tmp_812 <= 0;
      _tmp_813 <= 0;
      _tmp_814 <= 0;
      _tmp_815 <= 0;
      _tmp_816 <= 0;
      _tmp_817 <= 0;
      _tmp_818 <= 0;
      _tmp_819 <= 0;
      _tmp_820 <= 0;
      _tmp_821 <= 0;
      _tmp_822 <= 0;
      _tmp_823 <= 0;
      _tmp_824 <= 0;
      _tmp_825 <= 0;
      _tmp_826 <= 0;
      _tmp_827 <= 0;
      _tmp_828 <= 0;
      _tmp_829 <= 0;
      _tmp_830 <= 0;
      _tmp_831 <= 0;
      _tmp_832 <= 0;
      _tmp_833 <= 0;
      _tmp_834 <= 0;
      _tmp_835 <= 0;
      _tmp_836 <= 0;
      _tmp_837 <= 0;
      _tmp_838 <= 0;
      _tmp_839 <= 0;
      _tmp_840 <= 0;
      _tmp_841 <= 0;
      _tmp_842 <= 0;
      _tmp_843 <= 0;
      _tmp_844 <= 0;
      _tmp_845 <= 0;
      _tmp_846 <= 0;
      _tmp_847 <= 0;
      _tmp_848 <= 0;
      _tmp_849 <= 0;
      _tmp_850 <= 0;
      _tmp_851 <= 0;
      _tmp_852 <= 0;
      _tmp_853 <= 0;
      _tmp_854 <= 0;
      _tmp_855 <= 0;
      _tmp_856 <= 0;
      _tmp_857 <= 0;
      _tmp_858 <= 0;
      _tmp_859 <= 0;
      _tmp_860 <= 0;
      _tmp_861 <= 0;
      _tmp_862 <= 0;
      _tmp_863 <= 0;
      _tmp_864 <= 0;
      _tmp_865 <= 0;
      _tmp_866 <= 0;
      _tmp_867 <= 0;
      _tmp_868 <= 0;
      _tmp_869 <= 0;
      _tmp_870 <= 0;
      _tmp_871 <= 0;
      _tmp_872 <= 0;
      _tmp_873 <= 0;
      _tmp_874 <= 0;
      _tmp_875 <= 0;
      _tmp_876 <= 0;
      _tmp_877 <= 0;
      _tmp_878 <= 0;
      _tmp_879 <= 0;
      _tmp_880 <= 0;
      _tmp_881 <= 0;
      _tmp_882 <= 0;
      _tmp_883 <= 0;
      _tmp_884 <= 0;
      _tmp_885 <= 0;
      _tmp_886 <= 0;
      _tmp_887 <= 0;
      _tmp_888 <= 0;
      _tmp_889 <= 0;
      _tmp_890 <= 0;
      _tmp_891 <= 0;
      _tmp_892 <= 0;
      _tmp_893 <= 0;
      _tmp_894 <= 0;
      _tmp_895 <= 0;
      _tmp_896 <= 0;
      _tmp_897 <= 0;
      _tmp_898 <= 0;
      _tmp_899 <= 0;
      _tmp_900 <= 0;
      _tmp_901 <= 0;
      _tmp_902 <= 0;
      _tmp_903 <= 0;
      _tmp_904 <= 0;
      _tmp_905 <= 0;
      _tmp_906 <= 0;
      _tmp_907 <= 0;
      _tmp_908 <= 0;
      _tmp_909 <= 0;
      _tmp_910 <= 0;
      _tmp_911 <= 0;
      _tmp_912 <= 0;
      _tmp_913 <= 0;
      _tmp_914 <= 0;
      _tmp_915 <= 0;
      _tmp_916 <= 0;
      _tmp_917 <= 0;
      _tmp_918 <= 0;
      _tmp_919 <= 0;
      _stream_conv2d_25_busy_reg <= 0;
    end else begin
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_7_source_ram_renable <= 0;
        _stream_conv2d_25_source_7_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_7_idle <= _stream_conv2d_25_source_7_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_9_source_ram_renable <= 0;
        _stream_conv2d_25_source_9_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_9_idle <= _stream_conv2d_25_source_9_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_11_source_ram_renable <= 0;
        _stream_conv2d_25_source_11_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_11_idle <= _stream_conv2d_25_source_11_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_13_source_ram_renable <= 0;
        _stream_conv2d_25_source_13_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_13_idle <= _stream_conv2d_25_source_13_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_15_source_ram_renable <= 0;
        _stream_conv2d_25_source_15_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_15_idle <= _stream_conv2d_25_source_15_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_20_source_ram_renable <= 0;
        _stream_conv2d_25_source_20_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_20_idle <= _stream_conv2d_25_source_20_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_21_source_ram_renable <= 0;
        _stream_conv2d_25_source_21_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_21_idle <= _stream_conv2d_25_source_21_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_22_source_ram_renable <= 0;
        _stream_conv2d_25_source_22_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_22_idle <= _stream_conv2d_25_source_22_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_23_source_ram_renable <= 0;
        _stream_conv2d_25_source_23_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_23_idle <= _stream_conv2d_25_source_23_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_24_source_ram_renable <= 0;
        _stream_conv2d_25_source_24_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_24_idle <= _stream_conv2d_25_source_24_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_25_source_ram_renable <= 0;
        _stream_conv2d_25_source_25_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_25_idle <= _stream_conv2d_25_source_25_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_26_source_ram_renable <= 0;
        _stream_conv2d_25_source_26_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_26_idle <= _stream_conv2d_25_source_26_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_27_source_ram_renable <= 0;
        _stream_conv2d_25_source_27_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_27_idle <= _stream_conv2d_25_source_27_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_28_source_ram_renable <= 0;
        _stream_conv2d_25_source_28_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_28_idle <= _stream_conv2d_25_source_28_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_29_source_ram_renable <= 0;
        _stream_conv2d_25_source_29_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_29_idle <= _stream_conv2d_25_source_29_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_30_source_ram_renable <= 0;
        _stream_conv2d_25_source_30_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_30_idle <= _stream_conv2d_25_source_30_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_31_source_ram_renable <= 0;
        _stream_conv2d_25_source_31_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_31_idle <= _stream_conv2d_25_source_31_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_32_source_ram_renable <= 0;
        _stream_conv2d_25_source_32_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_32_idle <= _stream_conv2d_25_source_32_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_33_source_ram_renable <= 0;
        _stream_conv2d_25_source_33_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_33_idle <= _stream_conv2d_25_source_33_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_34_source_ram_renable <= 0;
        _stream_conv2d_25_source_34_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_34_idle <= _stream_conv2d_25_source_34_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_35_source_ram_renable <= 0;
        _stream_conv2d_25_source_35_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_35_idle <= _stream_conv2d_25_source_35_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_36_source_ram_renable <= 0;
        _stream_conv2d_25_source_36_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_36_idle <= _stream_conv2d_25_source_36_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_37_source_ram_renable <= 0;
        _stream_conv2d_25_source_37_source_fifo_deq <= 0;
      end 
      _stream_conv2d_25_source_37_idle <= _stream_conv2d_25_source_37_idle;
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_sink_50_sink_wenable <= 0;
        _stream_conv2d_25_sink_50_sink_fifo_enq <= 0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_sink_51_sink_wenable <= 0;
        _stream_conv2d_25_sink_51_sink_fifo_enq <= 0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_1 <= _stream_conv2d_25_stream_ivalid;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_2 <= __stream_conv2d_25_stream_ivalid_1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_3 <= __stream_conv2d_25_stream_ivalid_2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_4 <= __stream_conv2d_25_stream_ivalid_3;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_5 <= __stream_conv2d_25_stream_ivalid_4;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_6 <= __stream_conv2d_25_stream_ivalid_5;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_7 <= __stream_conv2d_25_stream_ivalid_6;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_8 <= __stream_conv2d_25_stream_ivalid_7;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_9 <= __stream_conv2d_25_stream_ivalid_8;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_10 <= __stream_conv2d_25_stream_ivalid_9;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_11 <= __stream_conv2d_25_stream_ivalid_10;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_12 <= __stream_conv2d_25_stream_ivalid_11;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_13 <= __stream_conv2d_25_stream_ivalid_12;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_14 <= __stream_conv2d_25_stream_ivalid_13;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_15 <= __stream_conv2d_25_stream_ivalid_14;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_16 <= __stream_conv2d_25_stream_ivalid_15;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_17 <= __stream_conv2d_25_stream_ivalid_16;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_18 <= __stream_conv2d_25_stream_ivalid_17;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_19 <= __stream_conv2d_25_stream_ivalid_18;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_20 <= __stream_conv2d_25_stream_ivalid_19;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_21 <= __stream_conv2d_25_stream_ivalid_20;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_22 <= __stream_conv2d_25_stream_ivalid_21;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_23 <= __stream_conv2d_25_stream_ivalid_22;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_24 <= __stream_conv2d_25_stream_ivalid_23;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_25 <= __stream_conv2d_25_stream_ivalid_24;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_26 <= __stream_conv2d_25_stream_ivalid_25;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_27 <= __stream_conv2d_25_stream_ivalid_26;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_28 <= __stream_conv2d_25_stream_ivalid_27;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_29 <= __stream_conv2d_25_stream_ivalid_28;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_30 <= __stream_conv2d_25_stream_ivalid_29;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_31 <= __stream_conv2d_25_stream_ivalid_30;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_32 <= __stream_conv2d_25_stream_ivalid_31;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_33 <= __stream_conv2d_25_stream_ivalid_32;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __stream_conv2d_25_stream_ivalid_34 <= __stream_conv2d_25_stream_ivalid_33;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_339 <= stream_conv2d_25_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_343 <= stream_conv2d_25_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_346 <= stream_conv2d_25_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_349 <= stream_conv2d_25_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_353 <= stream_conv2d_25_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_356 <= stream_conv2d_25_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_359 <= stream_conv2d_25_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_363 <= stream_conv2d_25_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_366 <= stream_conv2d_25_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_369 <= stream_conv2d_25_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_373 <= stream_conv2d_25_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_376 <= stream_conv2d_25_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_379 <= stream_conv2d_25_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_383 <= stream_conv2d_25_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_386 <= stream_conv2d_25_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_389 <= stream_conv2d_25_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_393 <= stream_conv2d_25_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_396 <= stream_conv2d_25_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_399 <= stream_conv2d_25_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_403 <= stream_conv2d_25_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_406 <= stream_conv2d_25_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_409 <= stream_conv2d_25_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_413 <= stream_conv2d_25_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_416 <= stream_conv2d_25_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_419 <= stream_conv2d_25_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_423 <= stream_conv2d_25_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_426 <= stream_conv2d_25_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_429 <= stream_conv2d_25_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_433 <= stream_conv2d_25_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_436 <= stream_conv2d_25_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_439 <= stream_conv2d_25_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_443 <= stream_conv2d_25_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_446 <= stream_conv2d_25_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_449 <= stream_conv2d_25_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_453 <= stream_conv2d_25_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_456 <= stream_conv2d_25_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_459 <= stream_conv2d_25_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_463 <= stream_conv2d_25_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_466 <= stream_conv2d_25_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_469 <= stream_conv2d_25_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_473 <= stream_conv2d_25_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_476 <= stream_conv2d_25_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_479 <= stream_conv2d_25_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_483 <= stream_conv2d_25_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_486 <= stream_conv2d_25_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_489 <= stream_conv2d_25_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_493 <= stream_conv2d_25_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_496 <= stream_conv2d_25_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_499 <= stream_conv2d_25_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_503 <= stream_conv2d_25_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_506 <= stream_conv2d_25_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_509 <= stream_conv2d_25_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_513 <= stream_conv2d_25_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _eq_data_516 <= stream_conv2d_25_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _plus_data_671 <= _cond_data_311 + stream_conv2d_25_parameter_16_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _plus_data_690 <= _cond_data_311 + stream_conv2d_25_parameter_16_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _plus_data_709 <= _cond_data_311 + stream_conv2d_25_parameter_16_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _plus_data_728 <= _cond_data_311 + stream_conv2d_25_parameter_16_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _plus_data_747 <= _cond_data_311 + stream_conv2d_25_parameter_16_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _plus_data_766 <= _cond_data_311 + stream_conv2d_25_parameter_16_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _plus_data_785 <= _cond_data_311 + stream_conv2d_25_parameter_16_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _plus_data_804 <= _cond_data_311 + stream_conv2d_25_parameter_16_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _plus_data_823 <= _cond_data_311 + stream_conv2d_25_parameter_16_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _plus_data_839 <= _cond_data_318 + stream_conv2d_25_parameter_17_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _plus_data_858 <= _cond_data_325 + stream_conv2d_25_parameter_18_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_946__variable_332 <= stream_conv2d_25_source_22_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_947__variable_331 <= stream_conv2d_25_source_21_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_948__variable_330 <= stream_conv2d_25_source_20_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_949__variable_335 <= stream_conv2d_25_source_25_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_950__variable_334 <= stream_conv2d_25_source_24_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_951__variable_333 <= stream_conv2d_25_source_23_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_952__variable_338 <= stream_conv2d_25_source_28_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_953__variable_337 <= stream_conv2d_25_source_27_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_954__variable_336 <= stream_conv2d_25_source_26_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_955_pointer_618 <= _pointer_data_618;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_956_reinterpretcast_609 <= _reinterpretcast_data_609;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_957_pointer_620 <= _pointer_data_620;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_958_reinterpretcast_610 <= _reinterpretcast_data_610;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_959_pointer_622 <= _pointer_data_622;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_960_reinterpretcast_611 <= _reinterpretcast_data_611;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_961_pointer_624 <= _pointer_data_624;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_962_reinterpretcast_612 <= _reinterpretcast_data_612;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_963_pointer_626 <= _pointer_data_626;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_964_reinterpretcast_613 <= _reinterpretcast_data_613;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_965_pointer_628 <= _pointer_data_628;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_966_reinterpretcast_614 <= _reinterpretcast_data_614;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_967_pointer_630 <= _pointer_data_630;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_968_reinterpretcast_615 <= _reinterpretcast_data_615;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_969_pointer_632 <= _pointer_data_632;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_970_reinterpretcast_616 <= _reinterpretcast_data_616;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_971_pointer_634 <= _pointer_data_634;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_972_reinterpretcast_617 <= _reinterpretcast_data_617;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_973__variable_281 <= stream_conv2d_25__reduce_reset_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_998__variable_276 <= stream_conv2d_25_parameter_0_data;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1011_cond_297 <= _cond_data_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1030_cond_304 <= _cond_data_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1069_eq_873 <= _eq_data_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_974__delay_973__variable_281 <= __delay_data_973__variable_281;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_986_plus_839 <= _plus_data_839;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_999__delay_998__variable_276 <= __delay_data_998__variable_276;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1012__delay_1011_cond_297 <= __delay_data_1011_cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1031__delay_1030_cond_304 <= __delay_data_1030_cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1050_plus_858 <= _plus_data_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1070__delay_1069_eq_873 <= __delay_data_1069_eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_975__delay_974__delay_973__variable_281 <= __delay_data_974__delay_973__variable_281;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_987__delay_986_plus_839 <= __delay_data_986_plus_839;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1000__delay_999__delay_998__variable_276 <= __delay_data_999__delay_998__variable_276;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1013__delay_1012__delay_1011_cond_297 <= __delay_data_1012__delay_1011_cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1032__delay_1031__delay_1030_cond_304 <= __delay_data_1031__delay_1030_cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1051__delay_1050_plus_858 <= __delay_data_1050_plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1071__delay_1070__delay_1069_eq_873 <= __delay_data_1070__delay_1069_eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_976__delay_975__delay_974____variable_281 <= __delay_data_975__delay_974__delay_973__variable_281;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_988__delay_987__delay_986_plus_839 <= __delay_data_987__delay_986_plus_839;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1001__delay_1000__delay_999____variable_276 <= __delay_data_1000__delay_999__delay_998__variable_276;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1014__delay_1013__delay_1012__delay_1011_cond_297 <= __delay_data_1013__delay_1012__delay_1011_cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1033__delay_1032__delay_1031__delay_1030_cond_304 <= __delay_data_1032__delay_1031__delay_1030_cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1052__delay_1051__delay_1050_plus_858 <= __delay_data_1051__delay_1050_plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1072__delay_1071__delay_1070__delay_1069_eq_873 <= __delay_data_1071__delay_1070__delay_1069_eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_977__delay_976__delay_975____variable_281 <= __delay_data_976__delay_975__delay_974____variable_281;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_989__delay_988__delay_987__delay_986_plus_839 <= __delay_data_988__delay_987__delay_986_plus_839;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1002__delay_1001__delay_1000____variable_276 <= __delay_data_1001__delay_1000__delay_999____variable_276;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1015__delay_1014__delay_1013__delay_1012___cond_297 <= __delay_data_1014__delay_1013__delay_1012__delay_1011_cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1034__delay_1033__delay_1032__delay_1031___cond_304 <= __delay_data_1033__delay_1032__delay_1031__delay_1030_cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1053__delay_1052__delay_1051__delay_1050_plus_858 <= __delay_data_1052__delay_1051__delay_1050_plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1073__delay_1072__delay_1071__delay_1070___eq_873 <= __delay_data_1072__delay_1071__delay_1070__delay_1069_eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_978__delay_977__delay_976____variable_281 <= __delay_data_977__delay_976__delay_975____variable_281;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_990__delay_989__delay_988__delay_987___plus_839 <= __delay_data_989__delay_988__delay_987__delay_986_plus_839;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1003__delay_1002__delay_1001____variable_276 <= __delay_data_1002__delay_1001__delay_1000____variable_276;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1016__delay_1015__delay_1014__delay_1013___cond_297 <= __delay_data_1015__delay_1014__delay_1013__delay_1012___cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1035__delay_1034__delay_1033__delay_1032___cond_304 <= __delay_data_1034__delay_1033__delay_1032__delay_1031___cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1054__delay_1053__delay_1052__delay_1051___plus_858 <= __delay_data_1053__delay_1052__delay_1051__delay_1050_plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1074__delay_1073__delay_1072__delay_1071___eq_873 <= __delay_data_1073__delay_1072__delay_1071__delay_1070___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_979__delay_978__delay_977____variable_281 <= __delay_data_978__delay_977__delay_976____variable_281;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_991__delay_990__delay_989__delay_988___plus_839 <= __delay_data_990__delay_989__delay_988__delay_987___plus_839;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1004__delay_1003__delay_1002____variable_276 <= __delay_data_1003__delay_1002__delay_1001____variable_276;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1017__delay_1016__delay_1015__delay_1014___cond_297 <= __delay_data_1016__delay_1015__delay_1014__delay_1013___cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1036__delay_1035__delay_1034__delay_1033___cond_304 <= __delay_data_1035__delay_1034__delay_1033__delay_1032___cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1055__delay_1054__delay_1053__delay_1052___plus_858 <= __delay_data_1054__delay_1053__delay_1052__delay_1051___plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1075__delay_1074__delay_1073__delay_1072___eq_873 <= __delay_data_1074__delay_1073__delay_1072__delay_1071___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_980__delay_979__delay_978____variable_281 <= __delay_data_979__delay_978__delay_977____variable_281;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_992__delay_991__delay_990__delay_989___plus_839 <= __delay_data_991__delay_990__delay_989__delay_988___plus_839;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1005__delay_1004__delay_1003____variable_276 <= __delay_data_1004__delay_1003__delay_1002____variable_276;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1018__delay_1017__delay_1016__delay_1015___cond_297 <= __delay_data_1017__delay_1016__delay_1015__delay_1014___cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1037__delay_1036__delay_1035__delay_1034___cond_304 <= __delay_data_1036__delay_1035__delay_1034__delay_1033___cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1056__delay_1055__delay_1054__delay_1053___plus_858 <= __delay_data_1055__delay_1054__delay_1053__delay_1052___plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1076__delay_1075__delay_1074__delay_1073___eq_873 <= __delay_data_1075__delay_1074__delay_1073__delay_1072___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_981__delay_980__delay_979____variable_281 <= __delay_data_980__delay_979__delay_978____variable_281;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_993__delay_992__delay_991__delay_990___plus_839 <= __delay_data_992__delay_991__delay_990__delay_989___plus_839;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1006__delay_1005__delay_1004____variable_276 <= __delay_data_1005__delay_1004__delay_1003____variable_276;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1019__delay_1018__delay_1017__delay_1016___cond_297 <= __delay_data_1018__delay_1017__delay_1016__delay_1015___cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1038__delay_1037__delay_1036__delay_1035___cond_304 <= __delay_data_1037__delay_1036__delay_1035__delay_1034___cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1057__delay_1056__delay_1055__delay_1054___plus_858 <= __delay_data_1056__delay_1055__delay_1054__delay_1053___plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1077__delay_1076__delay_1075__delay_1074___eq_873 <= __delay_data_1076__delay_1075__delay_1074__delay_1073___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_982__delay_981__delay_980____variable_281 <= __delay_data_981__delay_980__delay_979____variable_281;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_994__delay_993__delay_992__delay_991___plus_839 <= __delay_data_993__delay_992__delay_991__delay_990___plus_839;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1007__delay_1006__delay_1005____variable_276 <= __delay_data_1006__delay_1005__delay_1004____variable_276;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1020__delay_1019__delay_1018__delay_1017___cond_297 <= __delay_data_1019__delay_1018__delay_1017__delay_1016___cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1039__delay_1038__delay_1037__delay_1036___cond_304 <= __delay_data_1038__delay_1037__delay_1036__delay_1035___cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1058__delay_1057__delay_1056__delay_1055___plus_858 <= __delay_data_1057__delay_1056__delay_1055__delay_1054___plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1078__delay_1077__delay_1076__delay_1075___eq_873 <= __delay_data_1077__delay_1076__delay_1075__delay_1074___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_983__delay_982__delay_981____variable_281 <= __delay_data_982__delay_981__delay_980____variable_281;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_995__delay_994__delay_993__delay_992___plus_839 <= __delay_data_994__delay_993__delay_992__delay_991___plus_839;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1008__delay_1007__delay_1006____variable_276 <= __delay_data_1007__delay_1006__delay_1005____variable_276;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1021__delay_1020__delay_1019__delay_1018___cond_297 <= __delay_data_1020__delay_1019__delay_1018__delay_1017___cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1040__delay_1039__delay_1038__delay_1037___cond_304 <= __delay_data_1039__delay_1038__delay_1037__delay_1036___cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1059__delay_1058__delay_1057__delay_1056___plus_858 <= __delay_data_1058__delay_1057__delay_1056__delay_1055___plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1079__delay_1078__delay_1077__delay_1076___eq_873 <= __delay_data_1078__delay_1077__delay_1076__delay_1075___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_984__delay_983__delay_982____variable_281 <= __delay_data_983__delay_982__delay_981____variable_281;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_996__delay_995__delay_994__delay_993___plus_839 <= __delay_data_995__delay_994__delay_993__delay_992___plus_839;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1009__delay_1008__delay_1007____variable_276 <= __delay_data_1008__delay_1007__delay_1006____variable_276;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1022__delay_1021__delay_1020__delay_1019___cond_297 <= __delay_data_1021__delay_1020__delay_1019__delay_1018___cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1041__delay_1040__delay_1039__delay_1038___cond_304 <= __delay_data_1040__delay_1039__delay_1038__delay_1037___cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1060__delay_1059__delay_1058__delay_1057___plus_858 <= __delay_data_1059__delay_1058__delay_1057__delay_1056___plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1080__delay_1079__delay_1078__delay_1077___eq_873 <= __delay_data_1079__delay_1078__delay_1077__delay_1076___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_985__delay_984__delay_983____variable_281 <= __delay_data_984__delay_983__delay_982____variable_281;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_997__delay_996__delay_995__delay_994___plus_839 <= __delay_data_996__delay_995__delay_994__delay_993___plus_839;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1010__delay_1009__delay_1008____variable_276 <= __delay_data_1009__delay_1008__delay_1007____variable_276;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1023__delay_1022__delay_1021__delay_1020___cond_297 <= __delay_data_1022__delay_1021__delay_1020__delay_1019___cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1042__delay_1041__delay_1040__delay_1039___cond_304 <= __delay_data_1041__delay_1040__delay_1039__delay_1038___cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1061__delay_1060__delay_1059__delay_1058___plus_858 <= __delay_data_1060__delay_1059__delay_1058__delay_1057___plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1081__delay_1080__delay_1079__delay_1078___eq_873 <= __delay_data_1080__delay_1079__delay_1078__delay_1077___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1024__delay_1023__delay_1022__delay_1021___cond_297 <= __delay_data_1023__delay_1022__delay_1021__delay_1020___cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1043__delay_1042__delay_1041__delay_1040___cond_304 <= __delay_data_1042__delay_1041__delay_1040__delay_1039___cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1062__delay_1061__delay_1060__delay_1059___plus_858 <= __delay_data_1061__delay_1060__delay_1059__delay_1058___plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1082__delay_1081__delay_1080__delay_1079___eq_873 <= __delay_data_1081__delay_1080__delay_1079__delay_1078___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1025__delay_1024__delay_1023__delay_1022___cond_297 <= __delay_data_1024__delay_1023__delay_1022__delay_1021___cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1044__delay_1043__delay_1042__delay_1041___cond_304 <= __delay_data_1043__delay_1042__delay_1041__delay_1040___cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1063__delay_1062__delay_1061__delay_1060___plus_858 <= __delay_data_1062__delay_1061__delay_1060__delay_1059___plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1083__delay_1082__delay_1081__delay_1080___eq_873 <= __delay_data_1082__delay_1081__delay_1080__delay_1079___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1026__delay_1025__delay_1024__delay_1023___cond_297 <= __delay_data_1025__delay_1024__delay_1023__delay_1022___cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1045__delay_1044__delay_1043__delay_1042___cond_304 <= __delay_data_1044__delay_1043__delay_1042__delay_1041___cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1064__delay_1063__delay_1062__delay_1061___plus_858 <= __delay_data_1063__delay_1062__delay_1061__delay_1060___plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1084__delay_1083__delay_1082__delay_1081___eq_873 <= __delay_data_1083__delay_1082__delay_1081__delay_1080___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1027__delay_1026__delay_1025__delay_1024___cond_297 <= __delay_data_1026__delay_1025__delay_1024__delay_1023___cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1046__delay_1045__delay_1044__delay_1043___cond_304 <= __delay_data_1045__delay_1044__delay_1043__delay_1042___cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1065__delay_1064__delay_1063__delay_1062___plus_858 <= __delay_data_1064__delay_1063__delay_1062__delay_1061___plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1085__delay_1084__delay_1083__delay_1082___eq_873 <= __delay_data_1084__delay_1083__delay_1082__delay_1081___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1028__delay_1027__delay_1026__delay_1025___cond_297 <= __delay_data_1027__delay_1026__delay_1025__delay_1024___cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1047__delay_1046__delay_1045__delay_1044___cond_304 <= __delay_data_1046__delay_1045__delay_1044__delay_1043___cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1066__delay_1065__delay_1064__delay_1063___plus_858 <= __delay_data_1065__delay_1064__delay_1063__delay_1062___plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1086__delay_1085__delay_1084__delay_1083___eq_873 <= __delay_data_1085__delay_1084__delay_1083__delay_1082___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1029__delay_1028__delay_1027__delay_1026___cond_297 <= __delay_data_1028__delay_1027__delay_1026__delay_1025___cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1048__delay_1047__delay_1046__delay_1045___cond_304 <= __delay_data_1047__delay_1046__delay_1045__delay_1044___cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1067__delay_1066__delay_1065__delay_1064___plus_858 <= __delay_data_1066__delay_1065__delay_1064__delay_1063___plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1087__delay_1086__delay_1085__delay_1084___eq_873 <= __delay_data_1086__delay_1085__delay_1084__delay_1083___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _plus_data_842 <= __substreamoutput_data_840 + __delay_data_1029__delay_1028__delay_1027__delay_1026___cond_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1049__delay_1048__delay_1047__delay_1046___cond_304 <= __delay_data_1048__delay_1047__delay_1046__delay_1045___cond_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1068__delay_1067__delay_1066__delay_1065___plus_858 <= __delay_data_1067__delay_1066__delay_1065__delay_1064___plus_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1088__delay_1087__delay_1086__delay_1085___eq_873 <= __delay_data_1087__delay_1086__delay_1085__delay_1084___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1108__substreamoutput_841 <= __substreamoutput_data_841;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1089__delay_1088__delay_1087__delay_1086___eq_873 <= __delay_data_1088__delay_1087__delay_1086__delay_1085___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1109__delay_1108__substreamoutput_841 <= __delay_data_1108__substreamoutput_841;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1090__delay_1089__delay_1088__delay_1087___eq_873 <= __delay_data_1089__delay_1088__delay_1087__delay_1086___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1110__delay_1109__delay_1108__substreamoutput_841 <= __delay_data_1109__delay_1108__substreamoutput_841;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1091__delay_1090__delay_1089__delay_1088___eq_873 <= __delay_data_1090__delay_1089__delay_1088__delay_1087___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1111__delay_1110__delay_1109____substreamoutput_841 <= __delay_data_1110__delay_1109__delay_1108__substreamoutput_841;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1092__delay_1091__delay_1090__delay_1089___eq_873 <= __delay_data_1091__delay_1090__delay_1089__delay_1088___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1112__delay_1111__delay_1110____substreamoutput_841 <= __delay_data_1111__delay_1110__delay_1109____substreamoutput_841;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1093__delay_1092__delay_1091__delay_1090___eq_873 <= __delay_data_1092__delay_1091__delay_1090__delay_1089___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1113__delay_1112__delay_1111____substreamoutput_841 <= __delay_data_1112__delay_1111__delay_1110____substreamoutput_841;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1094__delay_1093__delay_1092__delay_1091___eq_873 <= __delay_data_1093__delay_1092__delay_1091__delay_1090___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1114__delay_1113__delay_1112____substreamoutput_841 <= __delay_data_1113__delay_1112__delay_1111____substreamoutput_841;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1095__delay_1094__delay_1093__delay_1092___eq_873 <= __delay_data_1094__delay_1093__delay_1092__delay_1091___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1115__delay_1114__delay_1113____substreamoutput_841 <= __delay_data_1114__delay_1113__delay_1112____substreamoutput_841;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1096__delay_1095__delay_1094__delay_1093___eq_873 <= __delay_data_1095__delay_1094__delay_1093__delay_1092___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1116__delay_1115__delay_1114____substreamoutput_841 <= __delay_data_1115__delay_1114__delay_1113____substreamoutput_841;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1097__delay_1096__delay_1095__delay_1094___eq_873 <= __delay_data_1096__delay_1095__delay_1094__delay_1093___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1117__delay_1116__delay_1115____substreamoutput_841 <= __delay_data_1116__delay_1115__delay_1114____substreamoutput_841;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _times_mul_odata_reg_860 <= _times_mul_odata_860;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _greaterthan_data_877 <= __substreamoutput_data_859 > 1'sd0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1098__delay_1097__delay_1096__delay_1095___eq_873 <= __delay_data_1097__delay_1096__delay_1095__delay_1094___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1104__substreamoutput_859 <= __substreamoutput_data_859;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1118__delay_1117__delay_1116____substreamoutput_841 <= __delay_data_1117__delay_1116__delay_1115____substreamoutput_841;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1099__delay_1098__delay_1097__delay_1096___eq_873 <= __delay_data_1098__delay_1097__delay_1096__delay_1095___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1101_greaterthan_877 <= _greaterthan_data_877;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1105__delay_1104__substreamoutput_859 <= __delay_data_1104__substreamoutput_859;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1119__delay_1118__delay_1117____substreamoutput_841 <= __delay_data_1118__delay_1117__delay_1116____substreamoutput_841;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1100__delay_1099__delay_1098__delay_1097___eq_873 <= __delay_data_1099__delay_1098__delay_1097__delay_1096___eq_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1102__delay_1101_greaterthan_877 <= __delay_data_1101_greaterthan_877;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1106__delay_1105__delay_1104__substreamoutput_859 <= __delay_data_1105__delay_1104__substreamoutput_859;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1120__delay_1119__delay_1118____substreamoutput_841 <= __delay_data_1119__delay_1118__delay_1117____substreamoutput_841;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _cond_data_875 <= (__delay_data_1100__delay_1099__delay_1098__delay_1097___eq_873)? _times_data_860 : _sra_data_870;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1103__delay_1102__delay_1101_greaterthan_877 <= __delay_data_1102__delay_1101_greaterthan_877;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1107__delay_1106__delay_1105____substreamoutput_859 <= __delay_data_1106__delay_1105__delay_1104__substreamoutput_859;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1121__delay_1120__delay_1119____substreamoutput_841 <= __delay_data_1120__delay_1119__delay_1118____substreamoutput_841;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _cond_data_878 <= (__delay_data_1103__delay_1102__delay_1101_greaterthan_877)? __delay_data_1107__delay_1106__delay_1105____substreamoutput_859 : _cond_data_875;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        __delay_data_1122__delay_1121__delay_1120____substreamoutput_841 <= __delay_data_1121__delay_1120__delay_1119____substreamoutput_841;
      end 
      if(_set_flag_218) begin
        _stream_conv2d_25_parameter_0_next_parameter_data <= cparam_conv2d_25_stream_reduce_size;
      end 
      if(_stream_conv2d_25_source_start) begin
        __variable_wdata_276 <= _stream_conv2d_25_parameter_0_next_parameter_data;
      end 
      if(_set_flag_219) begin
        _stream_conv2d_25_parameter_1_next_parameter_data <= conv2d_25_col_select;
      end 
      if(_stream_conv2d_25_source_start) begin
        __variable_wdata_277 <= _stream_conv2d_25_parameter_1_next_parameter_data;
      end 
      if(_set_flag_220) begin
        _stream_conv2d_25_parameter_2_next_parameter_data <= conv2d_25_row_select_buf;
      end 
      if(_stream_conv2d_25_source_start) begin
        __variable_wdata_278 <= _stream_conv2d_25_parameter_2_next_parameter_data;
      end 
      if(_set_flag_221) begin
        _stream_conv2d_25_parameter_3_next_parameter_data <= conv2d_25_stream_pad_masks;
      end 
      if(_stream_conv2d_25_source_start) begin
        __variable_wdata_279 <= _stream_conv2d_25_parameter_3_next_parameter_data;
      end 
      if(_set_flag_222) begin
        _stream_conv2d_25_parameter_4_next_parameter_data <= cparam_conv2d_25_stream_omit_mask;
      end 
      if(_stream_conv2d_25_source_start) begin
        __variable_wdata_280 <= _stream_conv2d_25_parameter_4_next_parameter_data;
      end 
      if(_set_flag_223) begin
        _stream_conv2d_25_parameter_6_next_parameter_data <= cparam_conv2d_25_bias_scala;
      end 
      if(_stream_conv2d_25_source_start) begin
        __variable_wdata_291 <= _stream_conv2d_25_parameter_6_next_parameter_data;
      end 
      if(_set_flag_224) begin
        _stream_conv2d_25_source_7_source_mode <= 5'b10;
        _stream_conv2d_25_source_7_source_offset <= (cparam_conv2d_25_bias_num == 1)? 0 : conv2d_25_och_count_buf;
      end 
      if(_set_flag_224) begin
        _source_stream_conv2d_25_source_7_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_7_pat_stride_0 <= 0;
      end 
      if(_set_flag_224) begin
        _source_stream_conv2d_25_source_7_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_7_pat_stride_1 <= (cparam_conv2d_25_bias_num == 1)? 0 : 1;
      end 
      if(_set_flag_224) begin
        _source_stream_conv2d_25_source_7_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_7_pat_stride_2 <= 0;
      end 
      if(_set_flag_224) begin
        _source_stream_conv2d_25_source_7_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_7_pat_stride_3 <= 0;
      end 
      if(_set_flag_224) begin
        _stream_conv2d_25_source_7_source_sel <= 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_7_source_offset_buf <= _stream_conv2d_25_source_7_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_count_0 <= _source_stream_conv2d_25_source_7_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_count_1 <= _source_stream_conv2d_25_source_7_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_count_2 <= _source_stream_conv2d_25_source_7_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_count_3 <= _source_stream_conv2d_25_source_7_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_size_buf_0 <= _source_stream_conv2d_25_source_7_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_size_buf_1 <= _source_stream_conv2d_25_source_7_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_size_buf_2 <= _source_stream_conv2d_25_source_7_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_size_buf_3 <= _source_stream_conv2d_25_source_7_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_stride_buf_0 <= _source_stream_conv2d_25_source_7_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_stride_buf_1 <= _source_stream_conv2d_25_source_7_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_stride_buf_2 <= _source_stream_conv2d_25_source_7_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_stride_buf_3 <= _source_stream_conv2d_25_source_7_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_292 <= _stream_conv2d_25_source_7_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_7_source_pat_fsm_0 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_7_idle <= 0;
        _stream_conv2d_25_source_7_source_ram_raddr <= _stream_conv2d_25_source_7_source_pat_all_offset;
        _stream_conv2d_25_source_7_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_7_source_pat_fsm_0 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_cur_offset_0 <= _source_stream_conv2d_25_source_7_pat_cur_offset_0 + _source_stream_conv2d_25_source_7_pat_stride_buf_0;
        _source_stream_conv2d_25_source_7_pat_count_0 <= _source_stream_conv2d_25_source_7_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_7_source_pat_fsm_0 == 1) && (_source_stream_conv2d_25_source_7_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_7_pat_count_0 <= _source_stream_conv2d_25_source_7_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_7_source_pat_fsm_0 == 1) && (_source_stream_conv2d_25_source_7_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_cur_offset_1 <= _source_stream_conv2d_25_source_7_pat_cur_offset_1 + _source_stream_conv2d_25_source_7_pat_stride_buf_1;
        _source_stream_conv2d_25_source_7_pat_count_1 <= _source_stream_conv2d_25_source_7_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_7_source_pat_fsm_0 == 1) && (_source_stream_conv2d_25_source_7_pat_count_0 == 0) && (_source_stream_conv2d_25_source_7_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_7_pat_count_1 <= _source_stream_conv2d_25_source_7_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_25_source_7_pat_count_0 == 0) && (_source_stream_conv2d_25_source_7_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_cur_offset_2 <= _source_stream_conv2d_25_source_7_pat_cur_offset_2 + _source_stream_conv2d_25_source_7_pat_stride_buf_2;
        _source_stream_conv2d_25_source_7_pat_count_2 <= _source_stream_conv2d_25_source_7_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_25_source_7_pat_count_0 == 0) && (_source_stream_conv2d_25_source_7_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_7_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_7_pat_count_2 <= _source_stream_conv2d_25_source_7_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_25_source_7_pat_count_0 == 0) && (_source_stream_conv2d_25_source_7_pat_count_1 == 0) && (_source_stream_conv2d_25_source_7_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_cur_offset_3 <= _source_stream_conv2d_25_source_7_pat_cur_offset_3 + _source_stream_conv2d_25_source_7_pat_stride_buf_3;
        _source_stream_conv2d_25_source_7_pat_count_3 <= _source_stream_conv2d_25_source_7_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_25_source_7_pat_count_0 == 0) && (_source_stream_conv2d_25_source_7_pat_count_1 == 0) && (_source_stream_conv2d_25_source_7_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_7_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_7_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_7_pat_count_3 <= _source_stream_conv2d_25_source_7_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_7_source_pat_fsm_0 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_7_source_ram_renable <= 0;
        _stream_conv2d_25_source_7_idle <= 1;
      end 
      if((_stream_conv2d_25_source_7_source_pat_fsm_0 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_7_source_ram_renable <= 0;
        _stream_conv2d_25_source_7_idle <= 1;
      end 
      if(_set_flag_227) begin
        _stream_conv2d_25_parameter_8_next_parameter_data <= cparam_conv2d_25_scale_scala;
      end 
      if(_stream_conv2d_25_source_start) begin
        __variable_wdata_298 <= _stream_conv2d_25_parameter_8_next_parameter_data;
      end 
      if(_set_flag_228) begin
        _stream_conv2d_25_source_9_source_mode <= 5'b10;
        _stream_conv2d_25_source_9_source_offset <= (cparam_conv2d_25_scale_num == 1)? 0 : conv2d_25_och_count_buf;
      end 
      if(_set_flag_228) begin
        _source_stream_conv2d_25_source_9_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_9_pat_stride_0 <= 0;
      end 
      if(_set_flag_228) begin
        _source_stream_conv2d_25_source_9_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_9_pat_stride_1 <= (cparam_conv2d_25_scale_num == 1)? 0 : 1;
      end 
      if(_set_flag_228) begin
        _source_stream_conv2d_25_source_9_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_9_pat_stride_2 <= 0;
      end 
      if(_set_flag_228) begin
        _source_stream_conv2d_25_source_9_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_9_pat_stride_3 <= 0;
      end 
      if(_set_flag_228) begin
        _stream_conv2d_25_source_9_source_sel <= 2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_9_source_offset_buf <= _stream_conv2d_25_source_9_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_count_0 <= _source_stream_conv2d_25_source_9_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_count_1 <= _source_stream_conv2d_25_source_9_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_count_2 <= _source_stream_conv2d_25_source_9_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_count_3 <= _source_stream_conv2d_25_source_9_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_size_buf_0 <= _source_stream_conv2d_25_source_9_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_size_buf_1 <= _source_stream_conv2d_25_source_9_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_size_buf_2 <= _source_stream_conv2d_25_source_9_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_size_buf_3 <= _source_stream_conv2d_25_source_9_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_stride_buf_0 <= _source_stream_conv2d_25_source_9_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_stride_buf_1 <= _source_stream_conv2d_25_source_9_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_stride_buf_2 <= _source_stream_conv2d_25_source_9_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_stride_buf_3 <= _source_stream_conv2d_25_source_9_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_299 <= _stream_conv2d_25_source_9_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_9_source_pat_fsm_1 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_9_idle <= 0;
        _stream_conv2d_25_source_9_source_ram_raddr <= _stream_conv2d_25_source_9_source_pat_all_offset;
        _stream_conv2d_25_source_9_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_9_source_pat_fsm_1 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_cur_offset_0 <= _source_stream_conv2d_25_source_9_pat_cur_offset_0 + _source_stream_conv2d_25_source_9_pat_stride_buf_0;
        _source_stream_conv2d_25_source_9_pat_count_0 <= _source_stream_conv2d_25_source_9_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_9_source_pat_fsm_1 == 1) && (_source_stream_conv2d_25_source_9_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_9_pat_count_0 <= _source_stream_conv2d_25_source_9_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_9_source_pat_fsm_1 == 1) && (_source_stream_conv2d_25_source_9_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_cur_offset_1 <= _source_stream_conv2d_25_source_9_pat_cur_offset_1 + _source_stream_conv2d_25_source_9_pat_stride_buf_1;
        _source_stream_conv2d_25_source_9_pat_count_1 <= _source_stream_conv2d_25_source_9_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_9_source_pat_fsm_1 == 1) && (_source_stream_conv2d_25_source_9_pat_count_0 == 0) && (_source_stream_conv2d_25_source_9_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_9_pat_count_1 <= _source_stream_conv2d_25_source_9_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_25_source_9_pat_count_0 == 0) && (_source_stream_conv2d_25_source_9_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_cur_offset_2 <= _source_stream_conv2d_25_source_9_pat_cur_offset_2 + _source_stream_conv2d_25_source_9_pat_stride_buf_2;
        _source_stream_conv2d_25_source_9_pat_count_2 <= _source_stream_conv2d_25_source_9_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_25_source_9_pat_count_0 == 0) && (_source_stream_conv2d_25_source_9_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_9_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_9_pat_count_2 <= _source_stream_conv2d_25_source_9_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_25_source_9_pat_count_0 == 0) && (_source_stream_conv2d_25_source_9_pat_count_1 == 0) && (_source_stream_conv2d_25_source_9_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_cur_offset_3 <= _source_stream_conv2d_25_source_9_pat_cur_offset_3 + _source_stream_conv2d_25_source_9_pat_stride_buf_3;
        _source_stream_conv2d_25_source_9_pat_count_3 <= _source_stream_conv2d_25_source_9_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_25_source_9_pat_count_0 == 0) && (_source_stream_conv2d_25_source_9_pat_count_1 == 0) && (_source_stream_conv2d_25_source_9_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_9_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_9_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_9_pat_count_3 <= _source_stream_conv2d_25_source_9_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_9_source_pat_fsm_1 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_9_source_ram_renable <= 0;
        _stream_conv2d_25_source_9_idle <= 1;
      end 
      if((_stream_conv2d_25_source_9_source_pat_fsm_1 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_9_source_ram_renable <= 0;
        _stream_conv2d_25_source_9_idle <= 1;
      end 
      if(_set_flag_231) begin
        _stream_conv2d_25_parameter_10_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_25_source_start) begin
        __variable_wdata_305 <= _stream_conv2d_25_parameter_10_next_parameter_data;
      end 
      if(_set_flag_232) begin
        _stream_conv2d_25_source_11_source_mode <= 5'b0;
        _stream_conv2d_25_source_11_source_empty_data <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_stream_oready && !(|(_stream_conv2d_25_source_11_source_mode & 5'b0))) begin
        _stream_conv2d_25_source_11_idle <= 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_stream_oready && !(|(_stream_conv2d_25_source_11_source_mode & 5'b0)) && _stream_conv2d_25_is_root) begin
        __variable_wdata_306 <= _stream_conv2d_25_source_11_source_empty_data;
      end 
      if(_set_flag_233) begin
        _stream_conv2d_25_parameter_12_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_25_source_start) begin
        __variable_wdata_312 <= _stream_conv2d_25_parameter_12_next_parameter_data;
      end 
      if(_set_flag_234) begin
        _stream_conv2d_25_source_13_source_mode <= 5'b0;
        _stream_conv2d_25_source_13_source_empty_data <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_stream_oready && !(|(_stream_conv2d_25_source_13_source_mode & 5'b0))) begin
        _stream_conv2d_25_source_13_idle <= 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_stream_oready && !(|(_stream_conv2d_25_source_13_source_mode & 5'b0)) && _stream_conv2d_25_is_root) begin
        __variable_wdata_313 <= _stream_conv2d_25_source_13_source_empty_data;
      end 
      if(_set_flag_235) begin
        _stream_conv2d_25_parameter_14_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_25_source_start) begin
        __variable_wdata_319 <= _stream_conv2d_25_parameter_14_next_parameter_data;
      end 
      if(_set_flag_236) begin
        _stream_conv2d_25_source_15_source_mode <= 5'b0;
        _stream_conv2d_25_source_15_source_empty_data <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_stream_oready && !(|(_stream_conv2d_25_source_15_source_mode & 5'b0))) begin
        _stream_conv2d_25_source_15_idle <= 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_stream_oready && !(|(_stream_conv2d_25_source_15_source_mode & 5'b0)) && _stream_conv2d_25_is_root) begin
        __variable_wdata_320 <= _stream_conv2d_25_source_15_source_empty_data;
      end 
      if(_set_flag_237) begin
        _stream_conv2d_25_parameter_16_next_parameter_data <= cparam_conv2d_25_cshamt_mul_value;
      end 
      if(_stream_conv2d_25_source_start) begin
        __variable_wdata_326 <= _stream_conv2d_25_parameter_16_next_parameter_data;
      end 
      if(_set_flag_238) begin
        _stream_conv2d_25_parameter_17_next_parameter_data <= cparam_conv2d_25_cshamt_sum_value;
      end 
      if(_stream_conv2d_25_source_start) begin
        __variable_wdata_327 <= _stream_conv2d_25_parameter_17_next_parameter_data;
      end 
      if(_set_flag_239) begin
        _stream_conv2d_25_parameter_18_next_parameter_data <= cparam_conv2d_25_cshamt_out_value;
      end 
      if(_stream_conv2d_25_source_start) begin
        __variable_wdata_328 <= _stream_conv2d_25_parameter_18_next_parameter_data;
      end 
      if(_set_flag_240) begin
        _stream_conv2d_25_parameter_19_next_parameter_data <= cparam_conv2d_25_act_func_index;
      end 
      if(_stream_conv2d_25_source_start) begin
        __variable_wdata_329 <= _stream_conv2d_25_parameter_19_next_parameter_data;
      end 
      if(_set_flag_241) begin
        _stream_conv2d_25_source_20_source_mode <= 5'b10;
        _stream_conv2d_25_source_20_source_offset <= conv2d_25_stream_act_local_0 + conv2d_25_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_241) begin
        _source_stream_conv2d_25_source_20_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_20_pat_stride_0 <= 1;
      end 
      if(_set_flag_241) begin
        _source_stream_conv2d_25_source_20_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_20_pat_stride_1 <= 0;
      end 
      if(_set_flag_241) begin
        _source_stream_conv2d_25_source_20_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_20_pat_stride_2 <= 0;
      end 
      if(_set_flag_241) begin
        _source_stream_conv2d_25_source_20_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_20_pat_stride_3 <= 0;
      end 
      if(_set_flag_241) begin
        _stream_conv2d_25_source_20_source_sel <= 3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_20_source_offset_buf <= _stream_conv2d_25_source_20_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_count_0 <= _source_stream_conv2d_25_source_20_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_count_1 <= _source_stream_conv2d_25_source_20_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_count_2 <= _source_stream_conv2d_25_source_20_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_count_3 <= _source_stream_conv2d_25_source_20_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_size_buf_0 <= _source_stream_conv2d_25_source_20_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_size_buf_1 <= _source_stream_conv2d_25_source_20_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_size_buf_2 <= _source_stream_conv2d_25_source_20_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_size_buf_3 <= _source_stream_conv2d_25_source_20_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_stride_buf_0 <= _source_stream_conv2d_25_source_20_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_stride_buf_1 <= _source_stream_conv2d_25_source_20_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_stride_buf_2 <= _source_stream_conv2d_25_source_20_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_stride_buf_3 <= _source_stream_conv2d_25_source_20_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_330 <= _stream_conv2d_25_source_20_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_20_source_pat_fsm_2 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_20_idle <= 0;
        _stream_conv2d_25_source_20_source_ram_raddr <= _stream_conv2d_25_source_20_source_pat_all_offset;
        _stream_conv2d_25_source_20_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_20_source_pat_fsm_2 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_cur_offset_0 <= _source_stream_conv2d_25_source_20_pat_cur_offset_0 + _source_stream_conv2d_25_source_20_pat_stride_buf_0;
        _source_stream_conv2d_25_source_20_pat_count_0 <= _source_stream_conv2d_25_source_20_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_20_source_pat_fsm_2 == 1) && (_source_stream_conv2d_25_source_20_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_20_pat_count_0 <= _source_stream_conv2d_25_source_20_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_20_source_pat_fsm_2 == 1) && (_source_stream_conv2d_25_source_20_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_cur_offset_1 <= _source_stream_conv2d_25_source_20_pat_cur_offset_1 + _source_stream_conv2d_25_source_20_pat_stride_buf_1;
        _source_stream_conv2d_25_source_20_pat_count_1 <= _source_stream_conv2d_25_source_20_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_20_source_pat_fsm_2 == 1) && (_source_stream_conv2d_25_source_20_pat_count_0 == 0) && (_source_stream_conv2d_25_source_20_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_20_pat_count_1 <= _source_stream_conv2d_25_source_20_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_25_source_20_pat_count_0 == 0) && (_source_stream_conv2d_25_source_20_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_cur_offset_2 <= _source_stream_conv2d_25_source_20_pat_cur_offset_2 + _source_stream_conv2d_25_source_20_pat_stride_buf_2;
        _source_stream_conv2d_25_source_20_pat_count_2 <= _source_stream_conv2d_25_source_20_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_25_source_20_pat_count_0 == 0) && (_source_stream_conv2d_25_source_20_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_20_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_20_pat_count_2 <= _source_stream_conv2d_25_source_20_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_25_source_20_pat_count_0 == 0) && (_source_stream_conv2d_25_source_20_pat_count_1 == 0) && (_source_stream_conv2d_25_source_20_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_cur_offset_3 <= _source_stream_conv2d_25_source_20_pat_cur_offset_3 + _source_stream_conv2d_25_source_20_pat_stride_buf_3;
        _source_stream_conv2d_25_source_20_pat_count_3 <= _source_stream_conv2d_25_source_20_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_25_source_20_pat_count_0 == 0) && (_source_stream_conv2d_25_source_20_pat_count_1 == 0) && (_source_stream_conv2d_25_source_20_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_20_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_20_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_20_pat_count_3 <= _source_stream_conv2d_25_source_20_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_20_source_pat_fsm_2 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_20_source_ram_renable <= 0;
        _stream_conv2d_25_source_20_idle <= 1;
      end 
      if((_stream_conv2d_25_source_20_source_pat_fsm_2 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_20_source_ram_renable <= 0;
        _stream_conv2d_25_source_20_idle <= 1;
      end 
      if(_set_flag_244) begin
        _stream_conv2d_25_source_21_source_mode <= 5'b10;
        _stream_conv2d_25_source_21_source_offset <= conv2d_25_stream_act_local_1 + conv2d_25_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_244) begin
        _source_stream_conv2d_25_source_21_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_21_pat_stride_0 <= 1;
      end 
      if(_set_flag_244) begin
        _source_stream_conv2d_25_source_21_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_21_pat_stride_1 <= 0;
      end 
      if(_set_flag_244) begin
        _source_stream_conv2d_25_source_21_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_21_pat_stride_2 <= 0;
      end 
      if(_set_flag_244) begin
        _source_stream_conv2d_25_source_21_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_21_pat_stride_3 <= 0;
      end 
      if(_set_flag_244) begin
        _stream_conv2d_25_source_21_source_sel <= 4;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_21_source_offset_buf <= _stream_conv2d_25_source_21_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_count_0 <= _source_stream_conv2d_25_source_21_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_count_1 <= _source_stream_conv2d_25_source_21_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_count_2 <= _source_stream_conv2d_25_source_21_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_count_3 <= _source_stream_conv2d_25_source_21_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_size_buf_0 <= _source_stream_conv2d_25_source_21_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_size_buf_1 <= _source_stream_conv2d_25_source_21_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_size_buf_2 <= _source_stream_conv2d_25_source_21_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_size_buf_3 <= _source_stream_conv2d_25_source_21_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_stride_buf_0 <= _source_stream_conv2d_25_source_21_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_stride_buf_1 <= _source_stream_conv2d_25_source_21_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_stride_buf_2 <= _source_stream_conv2d_25_source_21_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_stride_buf_3 <= _source_stream_conv2d_25_source_21_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_331 <= _stream_conv2d_25_source_21_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_21_source_pat_fsm_3 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_21_idle <= 0;
        _stream_conv2d_25_source_21_source_ram_raddr <= _stream_conv2d_25_source_21_source_pat_all_offset;
        _stream_conv2d_25_source_21_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_21_source_pat_fsm_3 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_cur_offset_0 <= _source_stream_conv2d_25_source_21_pat_cur_offset_0 + _source_stream_conv2d_25_source_21_pat_stride_buf_0;
        _source_stream_conv2d_25_source_21_pat_count_0 <= _source_stream_conv2d_25_source_21_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_21_source_pat_fsm_3 == 1) && (_source_stream_conv2d_25_source_21_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_21_pat_count_0 <= _source_stream_conv2d_25_source_21_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_21_source_pat_fsm_3 == 1) && (_source_stream_conv2d_25_source_21_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_cur_offset_1 <= _source_stream_conv2d_25_source_21_pat_cur_offset_1 + _source_stream_conv2d_25_source_21_pat_stride_buf_1;
        _source_stream_conv2d_25_source_21_pat_count_1 <= _source_stream_conv2d_25_source_21_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_21_source_pat_fsm_3 == 1) && (_source_stream_conv2d_25_source_21_pat_count_0 == 0) && (_source_stream_conv2d_25_source_21_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_21_pat_count_1 <= _source_stream_conv2d_25_source_21_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_25_source_21_pat_count_0 == 0) && (_source_stream_conv2d_25_source_21_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_cur_offset_2 <= _source_stream_conv2d_25_source_21_pat_cur_offset_2 + _source_stream_conv2d_25_source_21_pat_stride_buf_2;
        _source_stream_conv2d_25_source_21_pat_count_2 <= _source_stream_conv2d_25_source_21_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_25_source_21_pat_count_0 == 0) && (_source_stream_conv2d_25_source_21_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_21_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_21_pat_count_2 <= _source_stream_conv2d_25_source_21_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_25_source_21_pat_count_0 == 0) && (_source_stream_conv2d_25_source_21_pat_count_1 == 0) && (_source_stream_conv2d_25_source_21_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_cur_offset_3 <= _source_stream_conv2d_25_source_21_pat_cur_offset_3 + _source_stream_conv2d_25_source_21_pat_stride_buf_3;
        _source_stream_conv2d_25_source_21_pat_count_3 <= _source_stream_conv2d_25_source_21_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_25_source_21_pat_count_0 == 0) && (_source_stream_conv2d_25_source_21_pat_count_1 == 0) && (_source_stream_conv2d_25_source_21_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_21_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_21_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_21_pat_count_3 <= _source_stream_conv2d_25_source_21_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_21_source_pat_fsm_3 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_21_source_ram_renable <= 0;
        _stream_conv2d_25_source_21_idle <= 1;
      end 
      if((_stream_conv2d_25_source_21_source_pat_fsm_3 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_21_source_ram_renable <= 0;
        _stream_conv2d_25_source_21_idle <= 1;
      end 
      if(_set_flag_247) begin
        _stream_conv2d_25_source_22_source_mode <= 5'b10;
        _stream_conv2d_25_source_22_source_offset <= conv2d_25_stream_act_local_2 + conv2d_25_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_247) begin
        _source_stream_conv2d_25_source_22_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_22_pat_stride_0 <= 1;
      end 
      if(_set_flag_247) begin
        _source_stream_conv2d_25_source_22_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_22_pat_stride_1 <= 0;
      end 
      if(_set_flag_247) begin
        _source_stream_conv2d_25_source_22_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_22_pat_stride_2 <= 0;
      end 
      if(_set_flag_247) begin
        _source_stream_conv2d_25_source_22_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_22_pat_stride_3 <= 0;
      end 
      if(_set_flag_247) begin
        _stream_conv2d_25_source_22_source_sel <= 5;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_22_source_offset_buf <= _stream_conv2d_25_source_22_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_count_0 <= _source_stream_conv2d_25_source_22_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_count_1 <= _source_stream_conv2d_25_source_22_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_count_2 <= _source_stream_conv2d_25_source_22_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_count_3 <= _source_stream_conv2d_25_source_22_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_size_buf_0 <= _source_stream_conv2d_25_source_22_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_size_buf_1 <= _source_stream_conv2d_25_source_22_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_size_buf_2 <= _source_stream_conv2d_25_source_22_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_size_buf_3 <= _source_stream_conv2d_25_source_22_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_stride_buf_0 <= _source_stream_conv2d_25_source_22_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_stride_buf_1 <= _source_stream_conv2d_25_source_22_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_stride_buf_2 <= _source_stream_conv2d_25_source_22_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_stride_buf_3 <= _source_stream_conv2d_25_source_22_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_332 <= _stream_conv2d_25_source_22_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_22_source_pat_fsm_4 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_22_idle <= 0;
        _stream_conv2d_25_source_22_source_ram_raddr <= _stream_conv2d_25_source_22_source_pat_all_offset;
        _stream_conv2d_25_source_22_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_22_source_pat_fsm_4 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_cur_offset_0 <= _source_stream_conv2d_25_source_22_pat_cur_offset_0 + _source_stream_conv2d_25_source_22_pat_stride_buf_0;
        _source_stream_conv2d_25_source_22_pat_count_0 <= _source_stream_conv2d_25_source_22_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_22_source_pat_fsm_4 == 1) && (_source_stream_conv2d_25_source_22_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_22_pat_count_0 <= _source_stream_conv2d_25_source_22_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_22_source_pat_fsm_4 == 1) && (_source_stream_conv2d_25_source_22_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_cur_offset_1 <= _source_stream_conv2d_25_source_22_pat_cur_offset_1 + _source_stream_conv2d_25_source_22_pat_stride_buf_1;
        _source_stream_conv2d_25_source_22_pat_count_1 <= _source_stream_conv2d_25_source_22_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_22_source_pat_fsm_4 == 1) && (_source_stream_conv2d_25_source_22_pat_count_0 == 0) && (_source_stream_conv2d_25_source_22_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_22_pat_count_1 <= _source_stream_conv2d_25_source_22_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_25_source_22_pat_count_0 == 0) && (_source_stream_conv2d_25_source_22_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_cur_offset_2 <= _source_stream_conv2d_25_source_22_pat_cur_offset_2 + _source_stream_conv2d_25_source_22_pat_stride_buf_2;
        _source_stream_conv2d_25_source_22_pat_count_2 <= _source_stream_conv2d_25_source_22_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_25_source_22_pat_count_0 == 0) && (_source_stream_conv2d_25_source_22_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_22_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_22_pat_count_2 <= _source_stream_conv2d_25_source_22_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_25_source_22_pat_count_0 == 0) && (_source_stream_conv2d_25_source_22_pat_count_1 == 0) && (_source_stream_conv2d_25_source_22_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_cur_offset_3 <= _source_stream_conv2d_25_source_22_pat_cur_offset_3 + _source_stream_conv2d_25_source_22_pat_stride_buf_3;
        _source_stream_conv2d_25_source_22_pat_count_3 <= _source_stream_conv2d_25_source_22_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_25_source_22_pat_count_0 == 0) && (_source_stream_conv2d_25_source_22_pat_count_1 == 0) && (_source_stream_conv2d_25_source_22_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_22_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_22_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_22_pat_count_3 <= _source_stream_conv2d_25_source_22_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_22_source_pat_fsm_4 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_22_source_ram_renable <= 0;
        _stream_conv2d_25_source_22_idle <= 1;
      end 
      if((_stream_conv2d_25_source_22_source_pat_fsm_4 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_22_source_ram_renable <= 0;
        _stream_conv2d_25_source_22_idle <= 1;
      end 
      if(_set_flag_250) begin
        _stream_conv2d_25_source_23_source_mode <= 5'b10;
        _stream_conv2d_25_source_23_source_offset <= conv2d_25_stream_act_local_3 + conv2d_25_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_250) begin
        _source_stream_conv2d_25_source_23_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_23_pat_stride_0 <= 1;
      end 
      if(_set_flag_250) begin
        _source_stream_conv2d_25_source_23_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_23_pat_stride_1 <= 0;
      end 
      if(_set_flag_250) begin
        _source_stream_conv2d_25_source_23_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_23_pat_stride_2 <= 0;
      end 
      if(_set_flag_250) begin
        _source_stream_conv2d_25_source_23_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_23_pat_stride_3 <= 0;
      end 
      if(_set_flag_250) begin
        _stream_conv2d_25_source_23_source_sel <= 6;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_23_source_offset_buf <= _stream_conv2d_25_source_23_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_count_0 <= _source_stream_conv2d_25_source_23_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_count_1 <= _source_stream_conv2d_25_source_23_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_count_2 <= _source_stream_conv2d_25_source_23_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_count_3 <= _source_stream_conv2d_25_source_23_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_size_buf_0 <= _source_stream_conv2d_25_source_23_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_size_buf_1 <= _source_stream_conv2d_25_source_23_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_size_buf_2 <= _source_stream_conv2d_25_source_23_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_size_buf_3 <= _source_stream_conv2d_25_source_23_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_stride_buf_0 <= _source_stream_conv2d_25_source_23_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_stride_buf_1 <= _source_stream_conv2d_25_source_23_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_stride_buf_2 <= _source_stream_conv2d_25_source_23_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_stride_buf_3 <= _source_stream_conv2d_25_source_23_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_333 <= _stream_conv2d_25_source_23_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_23_source_pat_fsm_5 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_23_idle <= 0;
        _stream_conv2d_25_source_23_source_ram_raddr <= _stream_conv2d_25_source_23_source_pat_all_offset;
        _stream_conv2d_25_source_23_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_23_source_pat_fsm_5 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_cur_offset_0 <= _source_stream_conv2d_25_source_23_pat_cur_offset_0 + _source_stream_conv2d_25_source_23_pat_stride_buf_0;
        _source_stream_conv2d_25_source_23_pat_count_0 <= _source_stream_conv2d_25_source_23_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_23_source_pat_fsm_5 == 1) && (_source_stream_conv2d_25_source_23_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_23_pat_count_0 <= _source_stream_conv2d_25_source_23_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_23_source_pat_fsm_5 == 1) && (_source_stream_conv2d_25_source_23_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_cur_offset_1 <= _source_stream_conv2d_25_source_23_pat_cur_offset_1 + _source_stream_conv2d_25_source_23_pat_stride_buf_1;
        _source_stream_conv2d_25_source_23_pat_count_1 <= _source_stream_conv2d_25_source_23_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_23_source_pat_fsm_5 == 1) && (_source_stream_conv2d_25_source_23_pat_count_0 == 0) && (_source_stream_conv2d_25_source_23_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_23_pat_count_1 <= _source_stream_conv2d_25_source_23_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_25_source_23_pat_count_0 == 0) && (_source_stream_conv2d_25_source_23_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_cur_offset_2 <= _source_stream_conv2d_25_source_23_pat_cur_offset_2 + _source_stream_conv2d_25_source_23_pat_stride_buf_2;
        _source_stream_conv2d_25_source_23_pat_count_2 <= _source_stream_conv2d_25_source_23_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_25_source_23_pat_count_0 == 0) && (_source_stream_conv2d_25_source_23_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_23_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_23_pat_count_2 <= _source_stream_conv2d_25_source_23_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_25_source_23_pat_count_0 == 0) && (_source_stream_conv2d_25_source_23_pat_count_1 == 0) && (_source_stream_conv2d_25_source_23_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_cur_offset_3 <= _source_stream_conv2d_25_source_23_pat_cur_offset_3 + _source_stream_conv2d_25_source_23_pat_stride_buf_3;
        _source_stream_conv2d_25_source_23_pat_count_3 <= _source_stream_conv2d_25_source_23_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_25_source_23_pat_count_0 == 0) && (_source_stream_conv2d_25_source_23_pat_count_1 == 0) && (_source_stream_conv2d_25_source_23_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_23_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_23_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_23_pat_count_3 <= _source_stream_conv2d_25_source_23_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_23_source_pat_fsm_5 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_23_source_ram_renable <= 0;
        _stream_conv2d_25_source_23_idle <= 1;
      end 
      if((_stream_conv2d_25_source_23_source_pat_fsm_5 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_23_source_ram_renable <= 0;
        _stream_conv2d_25_source_23_idle <= 1;
      end 
      if(_set_flag_253) begin
        _stream_conv2d_25_source_24_source_mode <= 5'b10;
        _stream_conv2d_25_source_24_source_offset <= conv2d_25_stream_act_local_4 + conv2d_25_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_253) begin
        _source_stream_conv2d_25_source_24_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_24_pat_stride_0 <= 1;
      end 
      if(_set_flag_253) begin
        _source_stream_conv2d_25_source_24_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_24_pat_stride_1 <= 0;
      end 
      if(_set_flag_253) begin
        _source_stream_conv2d_25_source_24_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_24_pat_stride_2 <= 0;
      end 
      if(_set_flag_253) begin
        _source_stream_conv2d_25_source_24_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_24_pat_stride_3 <= 0;
      end 
      if(_set_flag_253) begin
        _stream_conv2d_25_source_24_source_sel <= 7;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_24_source_offset_buf <= _stream_conv2d_25_source_24_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_count_0 <= _source_stream_conv2d_25_source_24_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_count_1 <= _source_stream_conv2d_25_source_24_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_count_2 <= _source_stream_conv2d_25_source_24_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_count_3 <= _source_stream_conv2d_25_source_24_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_size_buf_0 <= _source_stream_conv2d_25_source_24_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_size_buf_1 <= _source_stream_conv2d_25_source_24_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_size_buf_2 <= _source_stream_conv2d_25_source_24_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_size_buf_3 <= _source_stream_conv2d_25_source_24_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_stride_buf_0 <= _source_stream_conv2d_25_source_24_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_stride_buf_1 <= _source_stream_conv2d_25_source_24_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_stride_buf_2 <= _source_stream_conv2d_25_source_24_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_stride_buf_3 <= _source_stream_conv2d_25_source_24_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_334 <= _stream_conv2d_25_source_24_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_24_source_pat_fsm_6 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_24_idle <= 0;
        _stream_conv2d_25_source_24_source_ram_raddr <= _stream_conv2d_25_source_24_source_pat_all_offset;
        _stream_conv2d_25_source_24_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_24_source_pat_fsm_6 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_cur_offset_0 <= _source_stream_conv2d_25_source_24_pat_cur_offset_0 + _source_stream_conv2d_25_source_24_pat_stride_buf_0;
        _source_stream_conv2d_25_source_24_pat_count_0 <= _source_stream_conv2d_25_source_24_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_24_source_pat_fsm_6 == 1) && (_source_stream_conv2d_25_source_24_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_24_pat_count_0 <= _source_stream_conv2d_25_source_24_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_24_source_pat_fsm_6 == 1) && (_source_stream_conv2d_25_source_24_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_cur_offset_1 <= _source_stream_conv2d_25_source_24_pat_cur_offset_1 + _source_stream_conv2d_25_source_24_pat_stride_buf_1;
        _source_stream_conv2d_25_source_24_pat_count_1 <= _source_stream_conv2d_25_source_24_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_24_source_pat_fsm_6 == 1) && (_source_stream_conv2d_25_source_24_pat_count_0 == 0) && (_source_stream_conv2d_25_source_24_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_24_pat_count_1 <= _source_stream_conv2d_25_source_24_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_25_source_24_pat_count_0 == 0) && (_source_stream_conv2d_25_source_24_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_cur_offset_2 <= _source_stream_conv2d_25_source_24_pat_cur_offset_2 + _source_stream_conv2d_25_source_24_pat_stride_buf_2;
        _source_stream_conv2d_25_source_24_pat_count_2 <= _source_stream_conv2d_25_source_24_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_25_source_24_pat_count_0 == 0) && (_source_stream_conv2d_25_source_24_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_24_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_24_pat_count_2 <= _source_stream_conv2d_25_source_24_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_25_source_24_pat_count_0 == 0) && (_source_stream_conv2d_25_source_24_pat_count_1 == 0) && (_source_stream_conv2d_25_source_24_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_cur_offset_3 <= _source_stream_conv2d_25_source_24_pat_cur_offset_3 + _source_stream_conv2d_25_source_24_pat_stride_buf_3;
        _source_stream_conv2d_25_source_24_pat_count_3 <= _source_stream_conv2d_25_source_24_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_25_source_24_pat_count_0 == 0) && (_source_stream_conv2d_25_source_24_pat_count_1 == 0) && (_source_stream_conv2d_25_source_24_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_24_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_24_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_24_pat_count_3 <= _source_stream_conv2d_25_source_24_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_24_source_pat_fsm_6 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_24_source_ram_renable <= 0;
        _stream_conv2d_25_source_24_idle <= 1;
      end 
      if((_stream_conv2d_25_source_24_source_pat_fsm_6 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_24_source_ram_renable <= 0;
        _stream_conv2d_25_source_24_idle <= 1;
      end 
      if(_set_flag_256) begin
        _stream_conv2d_25_source_25_source_mode <= 5'b10;
        _stream_conv2d_25_source_25_source_offset <= conv2d_25_stream_act_local_5 + conv2d_25_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_256) begin
        _source_stream_conv2d_25_source_25_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_25_pat_stride_0 <= 1;
      end 
      if(_set_flag_256) begin
        _source_stream_conv2d_25_source_25_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_25_pat_stride_1 <= 0;
      end 
      if(_set_flag_256) begin
        _source_stream_conv2d_25_source_25_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_25_pat_stride_2 <= 0;
      end 
      if(_set_flag_256) begin
        _source_stream_conv2d_25_source_25_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_25_pat_stride_3 <= 0;
      end 
      if(_set_flag_256) begin
        _stream_conv2d_25_source_25_source_sel <= 8;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_25_source_offset_buf <= _stream_conv2d_25_source_25_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_count_0 <= _source_stream_conv2d_25_source_25_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_count_1 <= _source_stream_conv2d_25_source_25_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_count_2 <= _source_stream_conv2d_25_source_25_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_count_3 <= _source_stream_conv2d_25_source_25_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_size_buf_0 <= _source_stream_conv2d_25_source_25_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_size_buf_1 <= _source_stream_conv2d_25_source_25_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_size_buf_2 <= _source_stream_conv2d_25_source_25_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_size_buf_3 <= _source_stream_conv2d_25_source_25_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_stride_buf_0 <= _source_stream_conv2d_25_source_25_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_stride_buf_1 <= _source_stream_conv2d_25_source_25_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_stride_buf_2 <= _source_stream_conv2d_25_source_25_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_stride_buf_3 <= _source_stream_conv2d_25_source_25_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_335 <= _stream_conv2d_25_source_25_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_25_source_pat_fsm_7 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_25_idle <= 0;
        _stream_conv2d_25_source_25_source_ram_raddr <= _stream_conv2d_25_source_25_source_pat_all_offset;
        _stream_conv2d_25_source_25_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_25_source_pat_fsm_7 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_cur_offset_0 <= _source_stream_conv2d_25_source_25_pat_cur_offset_0 + _source_stream_conv2d_25_source_25_pat_stride_buf_0;
        _source_stream_conv2d_25_source_25_pat_count_0 <= _source_stream_conv2d_25_source_25_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_25_source_pat_fsm_7 == 1) && (_source_stream_conv2d_25_source_25_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_25_pat_count_0 <= _source_stream_conv2d_25_source_25_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_25_source_pat_fsm_7 == 1) && (_source_stream_conv2d_25_source_25_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_cur_offset_1 <= _source_stream_conv2d_25_source_25_pat_cur_offset_1 + _source_stream_conv2d_25_source_25_pat_stride_buf_1;
        _source_stream_conv2d_25_source_25_pat_count_1 <= _source_stream_conv2d_25_source_25_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_25_source_pat_fsm_7 == 1) && (_source_stream_conv2d_25_source_25_pat_count_0 == 0) && (_source_stream_conv2d_25_source_25_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_25_pat_count_1 <= _source_stream_conv2d_25_source_25_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_25_source_25_pat_count_0 == 0) && (_source_stream_conv2d_25_source_25_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_cur_offset_2 <= _source_stream_conv2d_25_source_25_pat_cur_offset_2 + _source_stream_conv2d_25_source_25_pat_stride_buf_2;
        _source_stream_conv2d_25_source_25_pat_count_2 <= _source_stream_conv2d_25_source_25_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_25_source_25_pat_count_0 == 0) && (_source_stream_conv2d_25_source_25_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_25_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_25_pat_count_2 <= _source_stream_conv2d_25_source_25_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_25_source_25_pat_count_0 == 0) && (_source_stream_conv2d_25_source_25_pat_count_1 == 0) && (_source_stream_conv2d_25_source_25_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_cur_offset_3 <= _source_stream_conv2d_25_source_25_pat_cur_offset_3 + _source_stream_conv2d_25_source_25_pat_stride_buf_3;
        _source_stream_conv2d_25_source_25_pat_count_3 <= _source_stream_conv2d_25_source_25_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_25_source_25_pat_count_0 == 0) && (_source_stream_conv2d_25_source_25_pat_count_1 == 0) && (_source_stream_conv2d_25_source_25_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_25_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_25_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_25_pat_count_3 <= _source_stream_conv2d_25_source_25_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_25_source_pat_fsm_7 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_25_source_ram_renable <= 0;
        _stream_conv2d_25_source_25_idle <= 1;
      end 
      if((_stream_conv2d_25_source_25_source_pat_fsm_7 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_25_source_ram_renable <= 0;
        _stream_conv2d_25_source_25_idle <= 1;
      end 
      if(_set_flag_259) begin
        _stream_conv2d_25_source_26_source_mode <= 5'b10;
        _stream_conv2d_25_source_26_source_offset <= conv2d_25_stream_act_local_6 + conv2d_25_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_259) begin
        _source_stream_conv2d_25_source_26_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_26_pat_stride_0 <= 1;
      end 
      if(_set_flag_259) begin
        _source_stream_conv2d_25_source_26_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_26_pat_stride_1 <= 0;
      end 
      if(_set_flag_259) begin
        _source_stream_conv2d_25_source_26_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_26_pat_stride_2 <= 0;
      end 
      if(_set_flag_259) begin
        _source_stream_conv2d_25_source_26_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_26_pat_stride_3 <= 0;
      end 
      if(_set_flag_259) begin
        _stream_conv2d_25_source_26_source_sel <= 9;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_26_source_offset_buf <= _stream_conv2d_25_source_26_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_count_0 <= _source_stream_conv2d_25_source_26_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_count_1 <= _source_stream_conv2d_25_source_26_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_count_2 <= _source_stream_conv2d_25_source_26_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_count_3 <= _source_stream_conv2d_25_source_26_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_size_buf_0 <= _source_stream_conv2d_25_source_26_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_size_buf_1 <= _source_stream_conv2d_25_source_26_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_size_buf_2 <= _source_stream_conv2d_25_source_26_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_size_buf_3 <= _source_stream_conv2d_25_source_26_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_stride_buf_0 <= _source_stream_conv2d_25_source_26_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_stride_buf_1 <= _source_stream_conv2d_25_source_26_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_stride_buf_2 <= _source_stream_conv2d_25_source_26_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_stride_buf_3 <= _source_stream_conv2d_25_source_26_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_336 <= _stream_conv2d_25_source_26_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_26_source_pat_fsm_8 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_26_idle <= 0;
        _stream_conv2d_25_source_26_source_ram_raddr <= _stream_conv2d_25_source_26_source_pat_all_offset;
        _stream_conv2d_25_source_26_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_26_source_pat_fsm_8 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_cur_offset_0 <= _source_stream_conv2d_25_source_26_pat_cur_offset_0 + _source_stream_conv2d_25_source_26_pat_stride_buf_0;
        _source_stream_conv2d_25_source_26_pat_count_0 <= _source_stream_conv2d_25_source_26_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_26_source_pat_fsm_8 == 1) && (_source_stream_conv2d_25_source_26_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_26_pat_count_0 <= _source_stream_conv2d_25_source_26_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_26_source_pat_fsm_8 == 1) && (_source_stream_conv2d_25_source_26_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_cur_offset_1 <= _source_stream_conv2d_25_source_26_pat_cur_offset_1 + _source_stream_conv2d_25_source_26_pat_stride_buf_1;
        _source_stream_conv2d_25_source_26_pat_count_1 <= _source_stream_conv2d_25_source_26_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_26_source_pat_fsm_8 == 1) && (_source_stream_conv2d_25_source_26_pat_count_0 == 0) && (_source_stream_conv2d_25_source_26_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_26_pat_count_1 <= _source_stream_conv2d_25_source_26_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_25_source_26_pat_count_0 == 0) && (_source_stream_conv2d_25_source_26_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_cur_offset_2 <= _source_stream_conv2d_25_source_26_pat_cur_offset_2 + _source_stream_conv2d_25_source_26_pat_stride_buf_2;
        _source_stream_conv2d_25_source_26_pat_count_2 <= _source_stream_conv2d_25_source_26_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_25_source_26_pat_count_0 == 0) && (_source_stream_conv2d_25_source_26_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_26_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_26_pat_count_2 <= _source_stream_conv2d_25_source_26_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_25_source_26_pat_count_0 == 0) && (_source_stream_conv2d_25_source_26_pat_count_1 == 0) && (_source_stream_conv2d_25_source_26_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_cur_offset_3 <= _source_stream_conv2d_25_source_26_pat_cur_offset_3 + _source_stream_conv2d_25_source_26_pat_stride_buf_3;
        _source_stream_conv2d_25_source_26_pat_count_3 <= _source_stream_conv2d_25_source_26_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_25_source_26_pat_count_0 == 0) && (_source_stream_conv2d_25_source_26_pat_count_1 == 0) && (_source_stream_conv2d_25_source_26_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_26_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_26_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_26_pat_count_3 <= _source_stream_conv2d_25_source_26_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_26_source_pat_fsm_8 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_26_source_ram_renable <= 0;
        _stream_conv2d_25_source_26_idle <= 1;
      end 
      if((_stream_conv2d_25_source_26_source_pat_fsm_8 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_26_source_ram_renable <= 0;
        _stream_conv2d_25_source_26_idle <= 1;
      end 
      if(_set_flag_262) begin
        _stream_conv2d_25_source_27_source_mode <= 5'b10;
        _stream_conv2d_25_source_27_source_offset <= conv2d_25_stream_act_local_7 + conv2d_25_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_262) begin
        _source_stream_conv2d_25_source_27_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_27_pat_stride_0 <= 1;
      end 
      if(_set_flag_262) begin
        _source_stream_conv2d_25_source_27_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_27_pat_stride_1 <= 0;
      end 
      if(_set_flag_262) begin
        _source_stream_conv2d_25_source_27_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_27_pat_stride_2 <= 0;
      end 
      if(_set_flag_262) begin
        _source_stream_conv2d_25_source_27_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_27_pat_stride_3 <= 0;
      end 
      if(_set_flag_262) begin
        _stream_conv2d_25_source_27_source_sel <= 10;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_27_source_offset_buf <= _stream_conv2d_25_source_27_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_count_0 <= _source_stream_conv2d_25_source_27_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_count_1 <= _source_stream_conv2d_25_source_27_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_count_2 <= _source_stream_conv2d_25_source_27_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_count_3 <= _source_stream_conv2d_25_source_27_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_size_buf_0 <= _source_stream_conv2d_25_source_27_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_size_buf_1 <= _source_stream_conv2d_25_source_27_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_size_buf_2 <= _source_stream_conv2d_25_source_27_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_size_buf_3 <= _source_stream_conv2d_25_source_27_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_stride_buf_0 <= _source_stream_conv2d_25_source_27_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_stride_buf_1 <= _source_stream_conv2d_25_source_27_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_stride_buf_2 <= _source_stream_conv2d_25_source_27_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_stride_buf_3 <= _source_stream_conv2d_25_source_27_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_337 <= _stream_conv2d_25_source_27_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_27_source_pat_fsm_9 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_27_idle <= 0;
        _stream_conv2d_25_source_27_source_ram_raddr <= _stream_conv2d_25_source_27_source_pat_all_offset;
        _stream_conv2d_25_source_27_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_27_source_pat_fsm_9 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_cur_offset_0 <= _source_stream_conv2d_25_source_27_pat_cur_offset_0 + _source_stream_conv2d_25_source_27_pat_stride_buf_0;
        _source_stream_conv2d_25_source_27_pat_count_0 <= _source_stream_conv2d_25_source_27_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_27_source_pat_fsm_9 == 1) && (_source_stream_conv2d_25_source_27_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_27_pat_count_0 <= _source_stream_conv2d_25_source_27_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_27_source_pat_fsm_9 == 1) && (_source_stream_conv2d_25_source_27_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_cur_offset_1 <= _source_stream_conv2d_25_source_27_pat_cur_offset_1 + _source_stream_conv2d_25_source_27_pat_stride_buf_1;
        _source_stream_conv2d_25_source_27_pat_count_1 <= _source_stream_conv2d_25_source_27_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_27_source_pat_fsm_9 == 1) && (_source_stream_conv2d_25_source_27_pat_count_0 == 0) && (_source_stream_conv2d_25_source_27_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_27_pat_count_1 <= _source_stream_conv2d_25_source_27_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_25_source_27_pat_count_0 == 0) && (_source_stream_conv2d_25_source_27_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_cur_offset_2 <= _source_stream_conv2d_25_source_27_pat_cur_offset_2 + _source_stream_conv2d_25_source_27_pat_stride_buf_2;
        _source_stream_conv2d_25_source_27_pat_count_2 <= _source_stream_conv2d_25_source_27_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_25_source_27_pat_count_0 == 0) && (_source_stream_conv2d_25_source_27_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_27_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_27_pat_count_2 <= _source_stream_conv2d_25_source_27_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_25_source_27_pat_count_0 == 0) && (_source_stream_conv2d_25_source_27_pat_count_1 == 0) && (_source_stream_conv2d_25_source_27_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_cur_offset_3 <= _source_stream_conv2d_25_source_27_pat_cur_offset_3 + _source_stream_conv2d_25_source_27_pat_stride_buf_3;
        _source_stream_conv2d_25_source_27_pat_count_3 <= _source_stream_conv2d_25_source_27_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_25_source_27_pat_count_0 == 0) && (_source_stream_conv2d_25_source_27_pat_count_1 == 0) && (_source_stream_conv2d_25_source_27_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_27_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_27_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_27_pat_count_3 <= _source_stream_conv2d_25_source_27_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_27_source_pat_fsm_9 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_27_source_ram_renable <= 0;
        _stream_conv2d_25_source_27_idle <= 1;
      end 
      if((_stream_conv2d_25_source_27_source_pat_fsm_9 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_27_source_ram_renable <= 0;
        _stream_conv2d_25_source_27_idle <= 1;
      end 
      if(_set_flag_265) begin
        _stream_conv2d_25_source_28_source_mode <= 5'b10;
        _stream_conv2d_25_source_28_source_offset <= conv2d_25_stream_act_local_8 + conv2d_25_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_265) begin
        _source_stream_conv2d_25_source_28_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_28_pat_stride_0 <= 1;
      end 
      if(_set_flag_265) begin
        _source_stream_conv2d_25_source_28_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_28_pat_stride_1 <= 0;
      end 
      if(_set_flag_265) begin
        _source_stream_conv2d_25_source_28_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_28_pat_stride_2 <= 0;
      end 
      if(_set_flag_265) begin
        _source_stream_conv2d_25_source_28_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_28_pat_stride_3 <= 0;
      end 
      if(_set_flag_265) begin
        _stream_conv2d_25_source_28_source_sel <= 11;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_28_source_offset_buf <= _stream_conv2d_25_source_28_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_count_0 <= _source_stream_conv2d_25_source_28_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_count_1 <= _source_stream_conv2d_25_source_28_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_count_2 <= _source_stream_conv2d_25_source_28_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_count_3 <= _source_stream_conv2d_25_source_28_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_size_buf_0 <= _source_stream_conv2d_25_source_28_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_size_buf_1 <= _source_stream_conv2d_25_source_28_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_size_buf_2 <= _source_stream_conv2d_25_source_28_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_size_buf_3 <= _source_stream_conv2d_25_source_28_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_stride_buf_0 <= _source_stream_conv2d_25_source_28_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_stride_buf_1 <= _source_stream_conv2d_25_source_28_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_stride_buf_2 <= _source_stream_conv2d_25_source_28_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_stride_buf_3 <= _source_stream_conv2d_25_source_28_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_338 <= _stream_conv2d_25_source_28_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_28_source_pat_fsm_10 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_28_idle <= 0;
        _stream_conv2d_25_source_28_source_ram_raddr <= _stream_conv2d_25_source_28_source_pat_all_offset;
        _stream_conv2d_25_source_28_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_28_source_pat_fsm_10 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_cur_offset_0 <= _source_stream_conv2d_25_source_28_pat_cur_offset_0 + _source_stream_conv2d_25_source_28_pat_stride_buf_0;
        _source_stream_conv2d_25_source_28_pat_count_0 <= _source_stream_conv2d_25_source_28_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_28_source_pat_fsm_10 == 1) && (_source_stream_conv2d_25_source_28_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_28_pat_count_0 <= _source_stream_conv2d_25_source_28_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_28_source_pat_fsm_10 == 1) && (_source_stream_conv2d_25_source_28_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_cur_offset_1 <= _source_stream_conv2d_25_source_28_pat_cur_offset_1 + _source_stream_conv2d_25_source_28_pat_stride_buf_1;
        _source_stream_conv2d_25_source_28_pat_count_1 <= _source_stream_conv2d_25_source_28_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_28_source_pat_fsm_10 == 1) && (_source_stream_conv2d_25_source_28_pat_count_0 == 0) && (_source_stream_conv2d_25_source_28_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_28_pat_count_1 <= _source_stream_conv2d_25_source_28_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_25_source_28_pat_count_0 == 0) && (_source_stream_conv2d_25_source_28_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_cur_offset_2 <= _source_stream_conv2d_25_source_28_pat_cur_offset_2 + _source_stream_conv2d_25_source_28_pat_stride_buf_2;
        _source_stream_conv2d_25_source_28_pat_count_2 <= _source_stream_conv2d_25_source_28_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_25_source_28_pat_count_0 == 0) && (_source_stream_conv2d_25_source_28_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_28_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_28_pat_count_2 <= _source_stream_conv2d_25_source_28_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_25_source_28_pat_count_0 == 0) && (_source_stream_conv2d_25_source_28_pat_count_1 == 0) && (_source_stream_conv2d_25_source_28_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_cur_offset_3 <= _source_stream_conv2d_25_source_28_pat_cur_offset_3 + _source_stream_conv2d_25_source_28_pat_stride_buf_3;
        _source_stream_conv2d_25_source_28_pat_count_3 <= _source_stream_conv2d_25_source_28_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_25_source_28_pat_count_0 == 0) && (_source_stream_conv2d_25_source_28_pat_count_1 == 0) && (_source_stream_conv2d_25_source_28_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_28_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_28_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_28_pat_count_3 <= _source_stream_conv2d_25_source_28_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_28_source_pat_fsm_10 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_28_source_ram_renable <= 0;
        _stream_conv2d_25_source_28_idle <= 1;
      end 
      if((_stream_conv2d_25_source_28_source_pat_fsm_10 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_28_source_ram_renable <= 0;
        _stream_conv2d_25_source_28_idle <= 1;
      end 
      if(_set_flag_268) begin
        _stream_conv2d_25_source_29_source_mode <= 5'b10;
        _stream_conv2d_25_source_29_source_offset <= conv2d_25_filter_page_comp_offset_buf;
      end 
      if(_set_flag_268) begin
        _source_stream_conv2d_25_source_29_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_29_pat_stride_0 <= 1;
      end 
      if(_set_flag_268) begin
        _source_stream_conv2d_25_source_29_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_29_pat_stride_1 <= cparam_conv2d_25_stream_aligned_reduce_size;
      end 
      if(_set_flag_268) begin
        _source_stream_conv2d_25_source_29_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_29_pat_stride_2 <= 0;
      end 
      if(_set_flag_268) begin
        _source_stream_conv2d_25_source_29_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_29_pat_stride_3 <= 0;
      end 
      if(_set_flag_268) begin
        _stream_conv2d_25_source_29_source_sel <= 12;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_29_source_offset_buf <= _stream_conv2d_25_source_29_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_count_0 <= _source_stream_conv2d_25_source_29_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_count_1 <= _source_stream_conv2d_25_source_29_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_count_2 <= _source_stream_conv2d_25_source_29_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_count_3 <= _source_stream_conv2d_25_source_29_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_size_buf_0 <= _source_stream_conv2d_25_source_29_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_size_buf_1 <= _source_stream_conv2d_25_source_29_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_size_buf_2 <= _source_stream_conv2d_25_source_29_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_size_buf_3 <= _source_stream_conv2d_25_source_29_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_stride_buf_0 <= _source_stream_conv2d_25_source_29_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_stride_buf_1 <= _source_stream_conv2d_25_source_29_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_stride_buf_2 <= _source_stream_conv2d_25_source_29_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_stride_buf_3 <= _source_stream_conv2d_25_source_29_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_564 <= _stream_conv2d_25_source_29_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_29_source_pat_fsm_11 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_29_idle <= 0;
        _stream_conv2d_25_source_29_source_ram_raddr <= _stream_conv2d_25_source_29_source_pat_all_offset;
        _stream_conv2d_25_source_29_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_29_source_pat_fsm_11 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_cur_offset_0 <= _source_stream_conv2d_25_source_29_pat_cur_offset_0 + _source_stream_conv2d_25_source_29_pat_stride_buf_0;
        _source_stream_conv2d_25_source_29_pat_count_0 <= _source_stream_conv2d_25_source_29_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_29_source_pat_fsm_11 == 1) && (_source_stream_conv2d_25_source_29_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_29_pat_count_0 <= _source_stream_conv2d_25_source_29_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_29_source_pat_fsm_11 == 1) && (_source_stream_conv2d_25_source_29_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_cur_offset_1 <= _source_stream_conv2d_25_source_29_pat_cur_offset_1 + _source_stream_conv2d_25_source_29_pat_stride_buf_1;
        _source_stream_conv2d_25_source_29_pat_count_1 <= _source_stream_conv2d_25_source_29_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_29_source_pat_fsm_11 == 1) && (_source_stream_conv2d_25_source_29_pat_count_0 == 0) && (_source_stream_conv2d_25_source_29_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_29_pat_count_1 <= _source_stream_conv2d_25_source_29_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_25_source_29_pat_count_0 == 0) && (_source_stream_conv2d_25_source_29_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_cur_offset_2 <= _source_stream_conv2d_25_source_29_pat_cur_offset_2 + _source_stream_conv2d_25_source_29_pat_stride_buf_2;
        _source_stream_conv2d_25_source_29_pat_count_2 <= _source_stream_conv2d_25_source_29_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_25_source_29_pat_count_0 == 0) && (_source_stream_conv2d_25_source_29_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_29_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_29_pat_count_2 <= _source_stream_conv2d_25_source_29_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_25_source_29_pat_count_0 == 0) && (_source_stream_conv2d_25_source_29_pat_count_1 == 0) && (_source_stream_conv2d_25_source_29_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_cur_offset_3 <= _source_stream_conv2d_25_source_29_pat_cur_offset_3 + _source_stream_conv2d_25_source_29_pat_stride_buf_3;
        _source_stream_conv2d_25_source_29_pat_count_3 <= _source_stream_conv2d_25_source_29_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_25_source_29_pat_count_0 == 0) && (_source_stream_conv2d_25_source_29_pat_count_1 == 0) && (_source_stream_conv2d_25_source_29_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_29_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_29_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_29_pat_count_3 <= _source_stream_conv2d_25_source_29_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_29_source_pat_fsm_11 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_29_source_ram_renable <= 0;
        _stream_conv2d_25_source_29_idle <= 1;
      end 
      if((_stream_conv2d_25_source_29_source_pat_fsm_11 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_29_source_ram_renable <= 0;
        _stream_conv2d_25_source_29_idle <= 1;
      end 
      if(_set_flag_271) begin
        _stream_conv2d_25_source_30_source_mode <= 5'b10;
        _stream_conv2d_25_source_30_source_offset <= conv2d_25_filter_page_comp_offset_buf;
      end 
      if(_set_flag_271) begin
        _source_stream_conv2d_25_source_30_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_30_pat_stride_0 <= 1;
      end 
      if(_set_flag_271) begin
        _source_stream_conv2d_25_source_30_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_30_pat_stride_1 <= cparam_conv2d_25_stream_aligned_reduce_size;
      end 
      if(_set_flag_271) begin
        _source_stream_conv2d_25_source_30_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_30_pat_stride_2 <= 0;
      end 
      if(_set_flag_271) begin
        _source_stream_conv2d_25_source_30_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_30_pat_stride_3 <= 0;
      end 
      if(_set_flag_271) begin
        _stream_conv2d_25_source_30_source_sel <= 13;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_30_source_offset_buf <= _stream_conv2d_25_source_30_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_count_0 <= _source_stream_conv2d_25_source_30_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_count_1 <= _source_stream_conv2d_25_source_30_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_count_2 <= _source_stream_conv2d_25_source_30_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_count_3 <= _source_stream_conv2d_25_source_30_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_size_buf_0 <= _source_stream_conv2d_25_source_30_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_size_buf_1 <= _source_stream_conv2d_25_source_30_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_size_buf_2 <= _source_stream_conv2d_25_source_30_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_size_buf_3 <= _source_stream_conv2d_25_source_30_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_stride_buf_0 <= _source_stream_conv2d_25_source_30_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_stride_buf_1 <= _source_stream_conv2d_25_source_30_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_stride_buf_2 <= _source_stream_conv2d_25_source_30_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_stride_buf_3 <= _source_stream_conv2d_25_source_30_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_565 <= _stream_conv2d_25_source_30_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_30_source_pat_fsm_12 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_30_idle <= 0;
        _stream_conv2d_25_source_30_source_ram_raddr <= _stream_conv2d_25_source_30_source_pat_all_offset;
        _stream_conv2d_25_source_30_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_30_source_pat_fsm_12 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_cur_offset_0 <= _source_stream_conv2d_25_source_30_pat_cur_offset_0 + _source_stream_conv2d_25_source_30_pat_stride_buf_0;
        _source_stream_conv2d_25_source_30_pat_count_0 <= _source_stream_conv2d_25_source_30_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_30_source_pat_fsm_12 == 1) && (_source_stream_conv2d_25_source_30_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_30_pat_count_0 <= _source_stream_conv2d_25_source_30_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_30_source_pat_fsm_12 == 1) && (_source_stream_conv2d_25_source_30_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_cur_offset_1 <= _source_stream_conv2d_25_source_30_pat_cur_offset_1 + _source_stream_conv2d_25_source_30_pat_stride_buf_1;
        _source_stream_conv2d_25_source_30_pat_count_1 <= _source_stream_conv2d_25_source_30_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_30_source_pat_fsm_12 == 1) && (_source_stream_conv2d_25_source_30_pat_count_0 == 0) && (_source_stream_conv2d_25_source_30_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_30_pat_count_1 <= _source_stream_conv2d_25_source_30_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_25_source_30_pat_count_0 == 0) && (_source_stream_conv2d_25_source_30_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_cur_offset_2 <= _source_stream_conv2d_25_source_30_pat_cur_offset_2 + _source_stream_conv2d_25_source_30_pat_stride_buf_2;
        _source_stream_conv2d_25_source_30_pat_count_2 <= _source_stream_conv2d_25_source_30_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_25_source_30_pat_count_0 == 0) && (_source_stream_conv2d_25_source_30_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_30_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_30_pat_count_2 <= _source_stream_conv2d_25_source_30_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_25_source_30_pat_count_0 == 0) && (_source_stream_conv2d_25_source_30_pat_count_1 == 0) && (_source_stream_conv2d_25_source_30_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_cur_offset_3 <= _source_stream_conv2d_25_source_30_pat_cur_offset_3 + _source_stream_conv2d_25_source_30_pat_stride_buf_3;
        _source_stream_conv2d_25_source_30_pat_count_3 <= _source_stream_conv2d_25_source_30_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_25_source_30_pat_count_0 == 0) && (_source_stream_conv2d_25_source_30_pat_count_1 == 0) && (_source_stream_conv2d_25_source_30_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_30_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_30_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_30_pat_count_3 <= _source_stream_conv2d_25_source_30_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_30_source_pat_fsm_12 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_30_source_ram_renable <= 0;
        _stream_conv2d_25_source_30_idle <= 1;
      end 
      if((_stream_conv2d_25_source_30_source_pat_fsm_12 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_30_source_ram_renable <= 0;
        _stream_conv2d_25_source_30_idle <= 1;
      end 
      if(_set_flag_274) begin
        _stream_conv2d_25_source_31_source_mode <= 5'b10;
        _stream_conv2d_25_source_31_source_offset <= conv2d_25_filter_page_comp_offset_buf;
      end 
      if(_set_flag_274) begin
        _source_stream_conv2d_25_source_31_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_31_pat_stride_0 <= 1;
      end 
      if(_set_flag_274) begin
        _source_stream_conv2d_25_source_31_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_31_pat_stride_1 <= cparam_conv2d_25_stream_aligned_reduce_size;
      end 
      if(_set_flag_274) begin
        _source_stream_conv2d_25_source_31_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_31_pat_stride_2 <= 0;
      end 
      if(_set_flag_274) begin
        _source_stream_conv2d_25_source_31_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_31_pat_stride_3 <= 0;
      end 
      if(_set_flag_274) begin
        _stream_conv2d_25_source_31_source_sel <= 14;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_31_source_offset_buf <= _stream_conv2d_25_source_31_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_count_0 <= _source_stream_conv2d_25_source_31_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_count_1 <= _source_stream_conv2d_25_source_31_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_count_2 <= _source_stream_conv2d_25_source_31_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_count_3 <= _source_stream_conv2d_25_source_31_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_size_buf_0 <= _source_stream_conv2d_25_source_31_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_size_buf_1 <= _source_stream_conv2d_25_source_31_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_size_buf_2 <= _source_stream_conv2d_25_source_31_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_size_buf_3 <= _source_stream_conv2d_25_source_31_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_stride_buf_0 <= _source_stream_conv2d_25_source_31_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_stride_buf_1 <= _source_stream_conv2d_25_source_31_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_stride_buf_2 <= _source_stream_conv2d_25_source_31_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_stride_buf_3 <= _source_stream_conv2d_25_source_31_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_566 <= _stream_conv2d_25_source_31_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_31_source_pat_fsm_13 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_31_idle <= 0;
        _stream_conv2d_25_source_31_source_ram_raddr <= _stream_conv2d_25_source_31_source_pat_all_offset;
        _stream_conv2d_25_source_31_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_31_source_pat_fsm_13 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_cur_offset_0 <= _source_stream_conv2d_25_source_31_pat_cur_offset_0 + _source_stream_conv2d_25_source_31_pat_stride_buf_0;
        _source_stream_conv2d_25_source_31_pat_count_0 <= _source_stream_conv2d_25_source_31_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_31_source_pat_fsm_13 == 1) && (_source_stream_conv2d_25_source_31_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_31_pat_count_0 <= _source_stream_conv2d_25_source_31_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_31_source_pat_fsm_13 == 1) && (_source_stream_conv2d_25_source_31_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_cur_offset_1 <= _source_stream_conv2d_25_source_31_pat_cur_offset_1 + _source_stream_conv2d_25_source_31_pat_stride_buf_1;
        _source_stream_conv2d_25_source_31_pat_count_1 <= _source_stream_conv2d_25_source_31_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_31_source_pat_fsm_13 == 1) && (_source_stream_conv2d_25_source_31_pat_count_0 == 0) && (_source_stream_conv2d_25_source_31_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_31_pat_count_1 <= _source_stream_conv2d_25_source_31_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_25_source_31_pat_count_0 == 0) && (_source_stream_conv2d_25_source_31_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_cur_offset_2 <= _source_stream_conv2d_25_source_31_pat_cur_offset_2 + _source_stream_conv2d_25_source_31_pat_stride_buf_2;
        _source_stream_conv2d_25_source_31_pat_count_2 <= _source_stream_conv2d_25_source_31_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_25_source_31_pat_count_0 == 0) && (_source_stream_conv2d_25_source_31_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_31_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_31_pat_count_2 <= _source_stream_conv2d_25_source_31_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_25_source_31_pat_count_0 == 0) && (_source_stream_conv2d_25_source_31_pat_count_1 == 0) && (_source_stream_conv2d_25_source_31_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_cur_offset_3 <= _source_stream_conv2d_25_source_31_pat_cur_offset_3 + _source_stream_conv2d_25_source_31_pat_stride_buf_3;
        _source_stream_conv2d_25_source_31_pat_count_3 <= _source_stream_conv2d_25_source_31_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_25_source_31_pat_count_0 == 0) && (_source_stream_conv2d_25_source_31_pat_count_1 == 0) && (_source_stream_conv2d_25_source_31_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_31_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_31_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_31_pat_count_3 <= _source_stream_conv2d_25_source_31_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_31_source_pat_fsm_13 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_31_source_ram_renable <= 0;
        _stream_conv2d_25_source_31_idle <= 1;
      end 
      if((_stream_conv2d_25_source_31_source_pat_fsm_13 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_31_source_ram_renable <= 0;
        _stream_conv2d_25_source_31_idle <= 1;
      end 
      if(_set_flag_277) begin
        _stream_conv2d_25_source_32_source_mode <= 5'b10;
        _stream_conv2d_25_source_32_source_offset <= conv2d_25_filter_page_comp_offset_buf;
      end 
      if(_set_flag_277) begin
        _source_stream_conv2d_25_source_32_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_32_pat_stride_0 <= 1;
      end 
      if(_set_flag_277) begin
        _source_stream_conv2d_25_source_32_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_32_pat_stride_1 <= cparam_conv2d_25_stream_aligned_reduce_size;
      end 
      if(_set_flag_277) begin
        _source_stream_conv2d_25_source_32_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_32_pat_stride_2 <= 0;
      end 
      if(_set_flag_277) begin
        _source_stream_conv2d_25_source_32_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_32_pat_stride_3 <= 0;
      end 
      if(_set_flag_277) begin
        _stream_conv2d_25_source_32_source_sel <= 15;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_32_source_offset_buf <= _stream_conv2d_25_source_32_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_count_0 <= _source_stream_conv2d_25_source_32_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_count_1 <= _source_stream_conv2d_25_source_32_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_count_2 <= _source_stream_conv2d_25_source_32_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_count_3 <= _source_stream_conv2d_25_source_32_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_size_buf_0 <= _source_stream_conv2d_25_source_32_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_size_buf_1 <= _source_stream_conv2d_25_source_32_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_size_buf_2 <= _source_stream_conv2d_25_source_32_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_size_buf_3 <= _source_stream_conv2d_25_source_32_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_stride_buf_0 <= _source_stream_conv2d_25_source_32_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_stride_buf_1 <= _source_stream_conv2d_25_source_32_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_stride_buf_2 <= _source_stream_conv2d_25_source_32_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_stride_buf_3 <= _source_stream_conv2d_25_source_32_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_567 <= _stream_conv2d_25_source_32_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_32_source_pat_fsm_14 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_32_idle <= 0;
        _stream_conv2d_25_source_32_source_ram_raddr <= _stream_conv2d_25_source_32_source_pat_all_offset;
        _stream_conv2d_25_source_32_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_32_source_pat_fsm_14 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_cur_offset_0 <= _source_stream_conv2d_25_source_32_pat_cur_offset_0 + _source_stream_conv2d_25_source_32_pat_stride_buf_0;
        _source_stream_conv2d_25_source_32_pat_count_0 <= _source_stream_conv2d_25_source_32_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_32_source_pat_fsm_14 == 1) && (_source_stream_conv2d_25_source_32_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_32_pat_count_0 <= _source_stream_conv2d_25_source_32_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_32_source_pat_fsm_14 == 1) && (_source_stream_conv2d_25_source_32_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_cur_offset_1 <= _source_stream_conv2d_25_source_32_pat_cur_offset_1 + _source_stream_conv2d_25_source_32_pat_stride_buf_1;
        _source_stream_conv2d_25_source_32_pat_count_1 <= _source_stream_conv2d_25_source_32_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_32_source_pat_fsm_14 == 1) && (_source_stream_conv2d_25_source_32_pat_count_0 == 0) && (_source_stream_conv2d_25_source_32_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_32_pat_count_1 <= _source_stream_conv2d_25_source_32_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_25_source_32_pat_count_0 == 0) && (_source_stream_conv2d_25_source_32_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_cur_offset_2 <= _source_stream_conv2d_25_source_32_pat_cur_offset_2 + _source_stream_conv2d_25_source_32_pat_stride_buf_2;
        _source_stream_conv2d_25_source_32_pat_count_2 <= _source_stream_conv2d_25_source_32_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_25_source_32_pat_count_0 == 0) && (_source_stream_conv2d_25_source_32_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_32_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_32_pat_count_2 <= _source_stream_conv2d_25_source_32_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_25_source_32_pat_count_0 == 0) && (_source_stream_conv2d_25_source_32_pat_count_1 == 0) && (_source_stream_conv2d_25_source_32_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_cur_offset_3 <= _source_stream_conv2d_25_source_32_pat_cur_offset_3 + _source_stream_conv2d_25_source_32_pat_stride_buf_3;
        _source_stream_conv2d_25_source_32_pat_count_3 <= _source_stream_conv2d_25_source_32_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_25_source_32_pat_count_0 == 0) && (_source_stream_conv2d_25_source_32_pat_count_1 == 0) && (_source_stream_conv2d_25_source_32_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_32_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_32_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_32_pat_count_3 <= _source_stream_conv2d_25_source_32_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_32_source_pat_fsm_14 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_32_source_ram_renable <= 0;
        _stream_conv2d_25_source_32_idle <= 1;
      end 
      if((_stream_conv2d_25_source_32_source_pat_fsm_14 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_32_source_ram_renable <= 0;
        _stream_conv2d_25_source_32_idle <= 1;
      end 
      if(_set_flag_280) begin
        _stream_conv2d_25_source_33_source_mode <= 5'b10;
        _stream_conv2d_25_source_33_source_offset <= conv2d_25_filter_page_comp_offset_buf;
      end 
      if(_set_flag_280) begin
        _source_stream_conv2d_25_source_33_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_33_pat_stride_0 <= 1;
      end 
      if(_set_flag_280) begin
        _source_stream_conv2d_25_source_33_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_33_pat_stride_1 <= cparam_conv2d_25_stream_aligned_reduce_size;
      end 
      if(_set_flag_280) begin
        _source_stream_conv2d_25_source_33_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_33_pat_stride_2 <= 0;
      end 
      if(_set_flag_280) begin
        _source_stream_conv2d_25_source_33_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_33_pat_stride_3 <= 0;
      end 
      if(_set_flag_280) begin
        _stream_conv2d_25_source_33_source_sel <= 16;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_33_source_offset_buf <= _stream_conv2d_25_source_33_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_count_0 <= _source_stream_conv2d_25_source_33_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_count_1 <= _source_stream_conv2d_25_source_33_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_count_2 <= _source_stream_conv2d_25_source_33_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_count_3 <= _source_stream_conv2d_25_source_33_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_size_buf_0 <= _source_stream_conv2d_25_source_33_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_size_buf_1 <= _source_stream_conv2d_25_source_33_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_size_buf_2 <= _source_stream_conv2d_25_source_33_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_size_buf_3 <= _source_stream_conv2d_25_source_33_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_stride_buf_0 <= _source_stream_conv2d_25_source_33_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_stride_buf_1 <= _source_stream_conv2d_25_source_33_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_stride_buf_2 <= _source_stream_conv2d_25_source_33_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_stride_buf_3 <= _source_stream_conv2d_25_source_33_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_568 <= _stream_conv2d_25_source_33_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_33_source_pat_fsm_15 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_33_idle <= 0;
        _stream_conv2d_25_source_33_source_ram_raddr <= _stream_conv2d_25_source_33_source_pat_all_offset;
        _stream_conv2d_25_source_33_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_33_source_pat_fsm_15 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_cur_offset_0 <= _source_stream_conv2d_25_source_33_pat_cur_offset_0 + _source_stream_conv2d_25_source_33_pat_stride_buf_0;
        _source_stream_conv2d_25_source_33_pat_count_0 <= _source_stream_conv2d_25_source_33_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_33_source_pat_fsm_15 == 1) && (_source_stream_conv2d_25_source_33_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_33_pat_count_0 <= _source_stream_conv2d_25_source_33_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_33_source_pat_fsm_15 == 1) && (_source_stream_conv2d_25_source_33_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_cur_offset_1 <= _source_stream_conv2d_25_source_33_pat_cur_offset_1 + _source_stream_conv2d_25_source_33_pat_stride_buf_1;
        _source_stream_conv2d_25_source_33_pat_count_1 <= _source_stream_conv2d_25_source_33_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_33_source_pat_fsm_15 == 1) && (_source_stream_conv2d_25_source_33_pat_count_0 == 0) && (_source_stream_conv2d_25_source_33_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_33_pat_count_1 <= _source_stream_conv2d_25_source_33_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_25_source_33_pat_count_0 == 0) && (_source_stream_conv2d_25_source_33_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_cur_offset_2 <= _source_stream_conv2d_25_source_33_pat_cur_offset_2 + _source_stream_conv2d_25_source_33_pat_stride_buf_2;
        _source_stream_conv2d_25_source_33_pat_count_2 <= _source_stream_conv2d_25_source_33_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_25_source_33_pat_count_0 == 0) && (_source_stream_conv2d_25_source_33_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_33_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_33_pat_count_2 <= _source_stream_conv2d_25_source_33_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_25_source_33_pat_count_0 == 0) && (_source_stream_conv2d_25_source_33_pat_count_1 == 0) && (_source_stream_conv2d_25_source_33_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_cur_offset_3 <= _source_stream_conv2d_25_source_33_pat_cur_offset_3 + _source_stream_conv2d_25_source_33_pat_stride_buf_3;
        _source_stream_conv2d_25_source_33_pat_count_3 <= _source_stream_conv2d_25_source_33_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_25_source_33_pat_count_0 == 0) && (_source_stream_conv2d_25_source_33_pat_count_1 == 0) && (_source_stream_conv2d_25_source_33_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_33_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_33_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_33_pat_count_3 <= _source_stream_conv2d_25_source_33_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_33_source_pat_fsm_15 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_33_source_ram_renable <= 0;
        _stream_conv2d_25_source_33_idle <= 1;
      end 
      if((_stream_conv2d_25_source_33_source_pat_fsm_15 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_33_source_ram_renable <= 0;
        _stream_conv2d_25_source_33_idle <= 1;
      end 
      if(_set_flag_283) begin
        _stream_conv2d_25_source_34_source_mode <= 5'b10;
        _stream_conv2d_25_source_34_source_offset <= conv2d_25_filter_page_comp_offset_buf;
      end 
      if(_set_flag_283) begin
        _source_stream_conv2d_25_source_34_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_34_pat_stride_0 <= 1;
      end 
      if(_set_flag_283) begin
        _source_stream_conv2d_25_source_34_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_34_pat_stride_1 <= cparam_conv2d_25_stream_aligned_reduce_size;
      end 
      if(_set_flag_283) begin
        _source_stream_conv2d_25_source_34_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_34_pat_stride_2 <= 0;
      end 
      if(_set_flag_283) begin
        _source_stream_conv2d_25_source_34_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_34_pat_stride_3 <= 0;
      end 
      if(_set_flag_283) begin
        _stream_conv2d_25_source_34_source_sel <= 17;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_34_source_offset_buf <= _stream_conv2d_25_source_34_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_count_0 <= _source_stream_conv2d_25_source_34_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_count_1 <= _source_stream_conv2d_25_source_34_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_count_2 <= _source_stream_conv2d_25_source_34_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_count_3 <= _source_stream_conv2d_25_source_34_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_size_buf_0 <= _source_stream_conv2d_25_source_34_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_size_buf_1 <= _source_stream_conv2d_25_source_34_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_size_buf_2 <= _source_stream_conv2d_25_source_34_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_size_buf_3 <= _source_stream_conv2d_25_source_34_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_stride_buf_0 <= _source_stream_conv2d_25_source_34_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_stride_buf_1 <= _source_stream_conv2d_25_source_34_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_stride_buf_2 <= _source_stream_conv2d_25_source_34_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_stride_buf_3 <= _source_stream_conv2d_25_source_34_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_569 <= _stream_conv2d_25_source_34_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_34_source_pat_fsm_16 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_34_idle <= 0;
        _stream_conv2d_25_source_34_source_ram_raddr <= _stream_conv2d_25_source_34_source_pat_all_offset;
        _stream_conv2d_25_source_34_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_34_source_pat_fsm_16 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_cur_offset_0 <= _source_stream_conv2d_25_source_34_pat_cur_offset_0 + _source_stream_conv2d_25_source_34_pat_stride_buf_0;
        _source_stream_conv2d_25_source_34_pat_count_0 <= _source_stream_conv2d_25_source_34_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_34_source_pat_fsm_16 == 1) && (_source_stream_conv2d_25_source_34_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_34_pat_count_0 <= _source_stream_conv2d_25_source_34_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_34_source_pat_fsm_16 == 1) && (_source_stream_conv2d_25_source_34_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_cur_offset_1 <= _source_stream_conv2d_25_source_34_pat_cur_offset_1 + _source_stream_conv2d_25_source_34_pat_stride_buf_1;
        _source_stream_conv2d_25_source_34_pat_count_1 <= _source_stream_conv2d_25_source_34_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_34_source_pat_fsm_16 == 1) && (_source_stream_conv2d_25_source_34_pat_count_0 == 0) && (_source_stream_conv2d_25_source_34_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_34_pat_count_1 <= _source_stream_conv2d_25_source_34_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_25_source_34_pat_count_0 == 0) && (_source_stream_conv2d_25_source_34_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_cur_offset_2 <= _source_stream_conv2d_25_source_34_pat_cur_offset_2 + _source_stream_conv2d_25_source_34_pat_stride_buf_2;
        _source_stream_conv2d_25_source_34_pat_count_2 <= _source_stream_conv2d_25_source_34_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_25_source_34_pat_count_0 == 0) && (_source_stream_conv2d_25_source_34_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_34_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_34_pat_count_2 <= _source_stream_conv2d_25_source_34_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_25_source_34_pat_count_0 == 0) && (_source_stream_conv2d_25_source_34_pat_count_1 == 0) && (_source_stream_conv2d_25_source_34_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_cur_offset_3 <= _source_stream_conv2d_25_source_34_pat_cur_offset_3 + _source_stream_conv2d_25_source_34_pat_stride_buf_3;
        _source_stream_conv2d_25_source_34_pat_count_3 <= _source_stream_conv2d_25_source_34_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_25_source_34_pat_count_0 == 0) && (_source_stream_conv2d_25_source_34_pat_count_1 == 0) && (_source_stream_conv2d_25_source_34_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_34_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_34_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_34_pat_count_3 <= _source_stream_conv2d_25_source_34_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_34_source_pat_fsm_16 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_34_source_ram_renable <= 0;
        _stream_conv2d_25_source_34_idle <= 1;
      end 
      if((_stream_conv2d_25_source_34_source_pat_fsm_16 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_34_source_ram_renable <= 0;
        _stream_conv2d_25_source_34_idle <= 1;
      end 
      if(_set_flag_286) begin
        _stream_conv2d_25_source_35_source_mode <= 5'b10;
        _stream_conv2d_25_source_35_source_offset <= conv2d_25_filter_page_comp_offset_buf;
      end 
      if(_set_flag_286) begin
        _source_stream_conv2d_25_source_35_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_35_pat_stride_0 <= 1;
      end 
      if(_set_flag_286) begin
        _source_stream_conv2d_25_source_35_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_35_pat_stride_1 <= cparam_conv2d_25_stream_aligned_reduce_size;
      end 
      if(_set_flag_286) begin
        _source_stream_conv2d_25_source_35_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_35_pat_stride_2 <= 0;
      end 
      if(_set_flag_286) begin
        _source_stream_conv2d_25_source_35_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_35_pat_stride_3 <= 0;
      end 
      if(_set_flag_286) begin
        _stream_conv2d_25_source_35_source_sel <= 18;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_35_source_offset_buf <= _stream_conv2d_25_source_35_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_count_0 <= _source_stream_conv2d_25_source_35_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_count_1 <= _source_stream_conv2d_25_source_35_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_count_2 <= _source_stream_conv2d_25_source_35_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_count_3 <= _source_stream_conv2d_25_source_35_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_size_buf_0 <= _source_stream_conv2d_25_source_35_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_size_buf_1 <= _source_stream_conv2d_25_source_35_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_size_buf_2 <= _source_stream_conv2d_25_source_35_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_size_buf_3 <= _source_stream_conv2d_25_source_35_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_stride_buf_0 <= _source_stream_conv2d_25_source_35_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_stride_buf_1 <= _source_stream_conv2d_25_source_35_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_stride_buf_2 <= _source_stream_conv2d_25_source_35_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_stride_buf_3 <= _source_stream_conv2d_25_source_35_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_570 <= _stream_conv2d_25_source_35_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_35_source_pat_fsm_17 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_35_idle <= 0;
        _stream_conv2d_25_source_35_source_ram_raddr <= _stream_conv2d_25_source_35_source_pat_all_offset;
        _stream_conv2d_25_source_35_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_35_source_pat_fsm_17 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_cur_offset_0 <= _source_stream_conv2d_25_source_35_pat_cur_offset_0 + _source_stream_conv2d_25_source_35_pat_stride_buf_0;
        _source_stream_conv2d_25_source_35_pat_count_0 <= _source_stream_conv2d_25_source_35_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_35_source_pat_fsm_17 == 1) && (_source_stream_conv2d_25_source_35_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_35_pat_count_0 <= _source_stream_conv2d_25_source_35_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_35_source_pat_fsm_17 == 1) && (_source_stream_conv2d_25_source_35_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_cur_offset_1 <= _source_stream_conv2d_25_source_35_pat_cur_offset_1 + _source_stream_conv2d_25_source_35_pat_stride_buf_1;
        _source_stream_conv2d_25_source_35_pat_count_1 <= _source_stream_conv2d_25_source_35_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_35_source_pat_fsm_17 == 1) && (_source_stream_conv2d_25_source_35_pat_count_0 == 0) && (_source_stream_conv2d_25_source_35_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_35_pat_count_1 <= _source_stream_conv2d_25_source_35_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_25_source_35_pat_count_0 == 0) && (_source_stream_conv2d_25_source_35_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_cur_offset_2 <= _source_stream_conv2d_25_source_35_pat_cur_offset_2 + _source_stream_conv2d_25_source_35_pat_stride_buf_2;
        _source_stream_conv2d_25_source_35_pat_count_2 <= _source_stream_conv2d_25_source_35_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_25_source_35_pat_count_0 == 0) && (_source_stream_conv2d_25_source_35_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_35_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_35_pat_count_2 <= _source_stream_conv2d_25_source_35_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_25_source_35_pat_count_0 == 0) && (_source_stream_conv2d_25_source_35_pat_count_1 == 0) && (_source_stream_conv2d_25_source_35_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_cur_offset_3 <= _source_stream_conv2d_25_source_35_pat_cur_offset_3 + _source_stream_conv2d_25_source_35_pat_stride_buf_3;
        _source_stream_conv2d_25_source_35_pat_count_3 <= _source_stream_conv2d_25_source_35_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_25_source_35_pat_count_0 == 0) && (_source_stream_conv2d_25_source_35_pat_count_1 == 0) && (_source_stream_conv2d_25_source_35_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_35_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_35_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_35_pat_count_3 <= _source_stream_conv2d_25_source_35_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_35_source_pat_fsm_17 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_35_source_ram_renable <= 0;
        _stream_conv2d_25_source_35_idle <= 1;
      end 
      if((_stream_conv2d_25_source_35_source_pat_fsm_17 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_35_source_ram_renable <= 0;
        _stream_conv2d_25_source_35_idle <= 1;
      end 
      if(_set_flag_289) begin
        _stream_conv2d_25_source_36_source_mode <= 5'b10;
        _stream_conv2d_25_source_36_source_offset <= conv2d_25_filter_page_comp_offset_buf;
      end 
      if(_set_flag_289) begin
        _source_stream_conv2d_25_source_36_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_36_pat_stride_0 <= 1;
      end 
      if(_set_flag_289) begin
        _source_stream_conv2d_25_source_36_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_36_pat_stride_1 <= cparam_conv2d_25_stream_aligned_reduce_size;
      end 
      if(_set_flag_289) begin
        _source_stream_conv2d_25_source_36_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_36_pat_stride_2 <= 0;
      end 
      if(_set_flag_289) begin
        _source_stream_conv2d_25_source_36_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_36_pat_stride_3 <= 0;
      end 
      if(_set_flag_289) begin
        _stream_conv2d_25_source_36_source_sel <= 19;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_36_source_offset_buf <= _stream_conv2d_25_source_36_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_count_0 <= _source_stream_conv2d_25_source_36_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_count_1 <= _source_stream_conv2d_25_source_36_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_count_2 <= _source_stream_conv2d_25_source_36_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_count_3 <= _source_stream_conv2d_25_source_36_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_size_buf_0 <= _source_stream_conv2d_25_source_36_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_size_buf_1 <= _source_stream_conv2d_25_source_36_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_size_buf_2 <= _source_stream_conv2d_25_source_36_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_size_buf_3 <= _source_stream_conv2d_25_source_36_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_stride_buf_0 <= _source_stream_conv2d_25_source_36_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_stride_buf_1 <= _source_stream_conv2d_25_source_36_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_stride_buf_2 <= _source_stream_conv2d_25_source_36_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_stride_buf_3 <= _source_stream_conv2d_25_source_36_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_571 <= _stream_conv2d_25_source_36_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_36_source_pat_fsm_18 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_36_idle <= 0;
        _stream_conv2d_25_source_36_source_ram_raddr <= _stream_conv2d_25_source_36_source_pat_all_offset;
        _stream_conv2d_25_source_36_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_36_source_pat_fsm_18 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_cur_offset_0 <= _source_stream_conv2d_25_source_36_pat_cur_offset_0 + _source_stream_conv2d_25_source_36_pat_stride_buf_0;
        _source_stream_conv2d_25_source_36_pat_count_0 <= _source_stream_conv2d_25_source_36_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_36_source_pat_fsm_18 == 1) && (_source_stream_conv2d_25_source_36_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_36_pat_count_0 <= _source_stream_conv2d_25_source_36_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_36_source_pat_fsm_18 == 1) && (_source_stream_conv2d_25_source_36_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_cur_offset_1 <= _source_stream_conv2d_25_source_36_pat_cur_offset_1 + _source_stream_conv2d_25_source_36_pat_stride_buf_1;
        _source_stream_conv2d_25_source_36_pat_count_1 <= _source_stream_conv2d_25_source_36_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_36_source_pat_fsm_18 == 1) && (_source_stream_conv2d_25_source_36_pat_count_0 == 0) && (_source_stream_conv2d_25_source_36_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_36_pat_count_1 <= _source_stream_conv2d_25_source_36_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_25_source_36_pat_count_0 == 0) && (_source_stream_conv2d_25_source_36_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_cur_offset_2 <= _source_stream_conv2d_25_source_36_pat_cur_offset_2 + _source_stream_conv2d_25_source_36_pat_stride_buf_2;
        _source_stream_conv2d_25_source_36_pat_count_2 <= _source_stream_conv2d_25_source_36_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_25_source_36_pat_count_0 == 0) && (_source_stream_conv2d_25_source_36_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_36_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_36_pat_count_2 <= _source_stream_conv2d_25_source_36_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_25_source_36_pat_count_0 == 0) && (_source_stream_conv2d_25_source_36_pat_count_1 == 0) && (_source_stream_conv2d_25_source_36_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_cur_offset_3 <= _source_stream_conv2d_25_source_36_pat_cur_offset_3 + _source_stream_conv2d_25_source_36_pat_stride_buf_3;
        _source_stream_conv2d_25_source_36_pat_count_3 <= _source_stream_conv2d_25_source_36_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_25_source_36_pat_count_0 == 0) && (_source_stream_conv2d_25_source_36_pat_count_1 == 0) && (_source_stream_conv2d_25_source_36_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_36_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_36_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_36_pat_count_3 <= _source_stream_conv2d_25_source_36_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_36_source_pat_fsm_18 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_36_source_ram_renable <= 0;
        _stream_conv2d_25_source_36_idle <= 1;
      end 
      if((_stream_conv2d_25_source_36_source_pat_fsm_18 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_36_source_ram_renable <= 0;
        _stream_conv2d_25_source_36_idle <= 1;
      end 
      if(_set_flag_292) begin
        _stream_conv2d_25_source_37_source_mode <= 5'b10;
        _stream_conv2d_25_source_37_source_offset <= conv2d_25_filter_page_comp_offset_buf;
      end 
      if(_set_flag_292) begin
        _source_stream_conv2d_25_source_37_pat_size_0 <= cparam_conv2d_25_stream_reduce_size;
        _source_stream_conv2d_25_source_37_pat_stride_0 <= 1;
      end 
      if(_set_flag_292) begin
        _source_stream_conv2d_25_source_37_pat_size_1 <= conv2d_25_next_stream_num_ops;
        _source_stream_conv2d_25_source_37_pat_stride_1 <= cparam_conv2d_25_stream_aligned_reduce_size;
      end 
      if(_set_flag_292) begin
        _source_stream_conv2d_25_source_37_pat_size_2 <= 1;
        _source_stream_conv2d_25_source_37_pat_stride_2 <= 0;
      end 
      if(_set_flag_292) begin
        _source_stream_conv2d_25_source_37_pat_size_3 <= 1;
        _source_stream_conv2d_25_source_37_pat_stride_3 <= 0;
      end 
      if(_set_flag_292) begin
        _stream_conv2d_25_source_37_source_sel <= 20;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_37_source_offset_buf <= _stream_conv2d_25_source_37_source_offset;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_count_0 <= _source_stream_conv2d_25_source_37_pat_size_0 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_count_1 <= _source_stream_conv2d_25_source_37_pat_size_1 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_count_2 <= _source_stream_conv2d_25_source_37_pat_size_2 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_count_3 <= _source_stream_conv2d_25_source_37_pat_size_3 - 1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_size_buf_0 <= _source_stream_conv2d_25_source_37_pat_size_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_size_buf_1 <= _source_stream_conv2d_25_source_37_pat_size_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_size_buf_2 <= _source_stream_conv2d_25_source_37_pat_size_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_size_buf_3 <= _source_stream_conv2d_25_source_37_pat_size_3;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_stride_buf_0 <= _source_stream_conv2d_25_source_37_pat_stride_0;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_stride_buf_1 <= _source_stream_conv2d_25_source_37_pat_stride_1;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_stride_buf_2 <= _source_stream_conv2d_25_source_37_pat_stride_2;
      end 
      if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_stride_buf_3 <= _source_stream_conv2d_25_source_37_pat_stride_3;
      end 
      if(_stream_conv2d_25_stream_oready && _stream_conv2d_25_source_busy && _stream_conv2d_25_is_root) begin
        __variable_wdata_572 <= _stream_conv2d_25_source_37_source_ram_rdata;
      end 
      if((_stream_conv2d_25_source_37_source_pat_fsm_19 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_37_idle <= 0;
        _stream_conv2d_25_source_37_source_ram_raddr <= _stream_conv2d_25_source_37_source_pat_all_offset;
        _stream_conv2d_25_source_37_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_25_source_37_source_pat_fsm_19 == 1) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_cur_offset_0 <= _source_stream_conv2d_25_source_37_pat_cur_offset_0 + _source_stream_conv2d_25_source_37_pat_stride_buf_0;
        _source_stream_conv2d_25_source_37_pat_count_0 <= _source_stream_conv2d_25_source_37_pat_count_0 - 1;
      end 
      if((_stream_conv2d_25_source_37_source_pat_fsm_19 == 1) && (_source_stream_conv2d_25_source_37_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_25_source_37_pat_count_0 <= _source_stream_conv2d_25_source_37_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_25_source_37_source_pat_fsm_19 == 1) && (_source_stream_conv2d_25_source_37_pat_count_0 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_cur_offset_1 <= _source_stream_conv2d_25_source_37_pat_cur_offset_1 + _source_stream_conv2d_25_source_37_pat_stride_buf_1;
        _source_stream_conv2d_25_source_37_pat_count_1 <= _source_stream_conv2d_25_source_37_pat_count_1 - 1;
      end 
      if((_stream_conv2d_25_source_37_source_pat_fsm_19 == 1) && (_source_stream_conv2d_25_source_37_pat_count_0 == 0) && (_source_stream_conv2d_25_source_37_pat_count_1 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_25_source_37_pat_count_1 <= _source_stream_conv2d_25_source_37_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_25_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_25_source_37_pat_count_0 == 0) && (_source_stream_conv2d_25_source_37_pat_count_1 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_cur_offset_2 <= _source_stream_conv2d_25_source_37_pat_cur_offset_2 + _source_stream_conv2d_25_source_37_pat_stride_buf_2;
        _source_stream_conv2d_25_source_37_pat_count_2 <= _source_stream_conv2d_25_source_37_pat_count_2 - 1;
      end 
      if((_stream_conv2d_25_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_25_source_37_pat_count_0 == 0) && (_source_stream_conv2d_25_source_37_pat_count_1 == 0)) && (_source_stream_conv2d_25_source_37_pat_count_2 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_25_source_37_pat_count_2 <= _source_stream_conv2d_25_source_37_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_25_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_25_source_37_pat_count_0 == 0) && (_source_stream_conv2d_25_source_37_pat_count_1 == 0) && (_source_stream_conv2d_25_source_37_pat_count_2 == 0)) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_cur_offset_3 <= _source_stream_conv2d_25_source_37_pat_cur_offset_3 + _source_stream_conv2d_25_source_37_pat_stride_buf_3;
        _source_stream_conv2d_25_source_37_pat_count_3 <= _source_stream_conv2d_25_source_37_pat_count_3 - 1;
      end 
      if((_stream_conv2d_25_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_25_source_37_pat_count_0 == 0) && (_source_stream_conv2d_25_source_37_pat_count_1 == 0) && (_source_stream_conv2d_25_source_37_pat_count_2 == 0)) && (_source_stream_conv2d_25_source_37_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
        _source_stream_conv2d_25_source_37_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_25_source_37_pat_count_3 <= _source_stream_conv2d_25_source_37_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_25_source_37_source_pat_fsm_19 == 1) && _stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_37_source_ram_renable <= 0;
        _stream_conv2d_25_source_37_idle <= 1;
      end 
      if((_stream_conv2d_25_source_37_source_pat_fsm_19 == 2) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_source_37_source_ram_renable <= 0;
        _stream_conv2d_25_source_37_idle <= 1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_296 <= _set_flag_295;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_297 <= _tmp_296;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_298 <= _tmp_297;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_299 <= _tmp_298;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_300 <= _tmp_299;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_301 <= _tmp_300;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_302 <= _tmp_301;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_303 <= _tmp_302;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_304 <= _tmp_303;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_305 <= _tmp_304;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_306 <= _tmp_305;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_307 <= _tmp_306;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_308 <= _tmp_307;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_309 <= _tmp_308;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_310 <= _tmp_309;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_311 <= _tmp_310;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_312 <= _tmp_311;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_313 <= _tmp_312;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_314 <= _tmp_313;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_315 <= _tmp_314;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_316 <= _tmp_315;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_317 <= _tmp_316;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_318 <= _tmp_317;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_319 <= _tmp_318;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_320 <= _tmp_319;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_321 <= _tmp_320;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_322 <= _tmp_321;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_323 <= _tmp_322;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_324 <= _tmp_323;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_325 <= _tmp_324;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_326 <= _tmp_325;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_327 <= _tmp_326;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_328 <= _tmp_327;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_329 <= _tmp_328;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_330 <= _tmp_329;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_331 <= _tmp_330;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_334 <= _tmp_333;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_335 <= _tmp_334;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_336 <= _tmp_335;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_337 <= _tmp_336;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_338 <= _tmp_337;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_339 <= _tmp_338;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_340 <= _tmp_339;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_341 <= _tmp_340;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_342 <= _tmp_341;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_343 <= _tmp_342;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_344 <= _tmp_343;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_345 <= _tmp_344;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_346 <= _tmp_345;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_347 <= _tmp_346;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_348 <= _tmp_347;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_349 <= _tmp_348;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_350 <= _tmp_349;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_351 <= _tmp_350;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_352 <= _tmp_351;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_353 <= _tmp_352;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_354 <= _tmp_353;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_355 <= _tmp_354;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_356 <= _tmp_355;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_357 <= _tmp_356;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_358 <= _tmp_357;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_359 <= _tmp_358;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_360 <= _tmp_359;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_361 <= _tmp_360;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_362 <= _tmp_361;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_363 <= _tmp_362;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_364 <= _tmp_363;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_365 <= _tmp_364;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_366 <= _tmp_365;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_367 <= _tmp_366;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_368 <= _tmp_367;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_369 <= _tmp_368;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_370 <= conv2d_25_next_stream_num_ops;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_371 <= _tmp_370;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_372 <= _tmp_371;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_373 <= _tmp_372;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_374 <= _tmp_373;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_375 <= _tmp_374;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_376 <= _tmp_375;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_377 <= _tmp_376;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_378 <= _tmp_377;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_379 <= _tmp_378;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_380 <= _tmp_379;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_381 <= _tmp_380;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_382 <= _tmp_381;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_383 <= _tmp_382;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_384 <= _tmp_383;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_385 <= _tmp_384;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_386 <= _tmp_385;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_387 <= _tmp_386;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_388 <= _tmp_387;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_389 <= _tmp_388;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_390 <= _tmp_389;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_391 <= _tmp_390;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_392 <= _tmp_391;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_393 <= _tmp_392;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_394 <= _tmp_393;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_395 <= _tmp_394;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_396 <= _tmp_395;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_397 <= _tmp_396;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_398 <= _tmp_397;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_399 <= _tmp_398;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_400 <= _tmp_399;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_401 <= _tmp_400;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_402 <= _tmp_401;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_403 <= _tmp_402;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_404 <= _tmp_403;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_405 <= _tmp_404;
      end 
      if(_tmp_331) begin
        _stream_conv2d_25_sink_50_sink_mode <= 5'b1;
        _stream_conv2d_25_sink_50_sink_offset <= _tmp_369;
        _stream_conv2d_25_sink_50_sink_size <= _tmp_405;
        _stream_conv2d_25_sink_50_sink_stride <= 1;
      end 
      if(_tmp_331) begin
        _stream_conv2d_25_sink_50_sink_sel <= 21;
      end 
      if(_stream_conv2d_25_sink_start && _stream_conv2d_25_sink_50_sink_mode & 5'b1 && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_sink_50_sink_offset_buf <= _stream_conv2d_25_sink_50_sink_offset;
        _stream_conv2d_25_sink_50_sink_size_buf <= _stream_conv2d_25_sink_50_sink_size;
        _stream_conv2d_25_sink_50_sink_stride_buf <= _stream_conv2d_25_sink_50_sink_stride;
      end 
      if((_stream_conv2d_25_sink_50_sink_fsm_20 == 1) && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_sink_50_sink_waddr <= _stream_conv2d_25_sink_50_sink_offset_buf - _stream_conv2d_25_sink_50_sink_stride_buf;
        _stream_conv2d_25_sink_50_sink_count <= _stream_conv2d_25_sink_50_sink_size_buf;
      end 
      if((_stream_conv2d_25_sink_50_sink_fsm_20 == 2) && stream_conv2d_25_sink_51_data && _stream_conv2d_25_stream_oready) begin
        _stream_conv2d_25_sink_50_sink_waddr <= _stream_conv2d_25_sink_50_sink_waddr + _stream_conv2d_25_sink_50_sink_stride_buf;
        _stream_conv2d_25_sink_50_sink_wdata <= stream_conv2d_25_sink_50_data;
        _stream_conv2d_25_sink_50_sink_wenable <= 1;
        _stream_conv2d_25_sink_50_sink_count <= _stream_conv2d_25_sink_50_sink_count - 1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_795 <= _stream_conv2d_25_source_start;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_796 <= _tmp_795;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_797 <= _tmp_796;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_798 <= _stream_conv2d_25_source_start;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_799 <= _tmp_798;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_800 <= _tmp_799;
      end 
      if(_stream_conv2d_25_stream_oready && _tmp_800) begin
        __variable_wdata_281 <= 1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_801 <= _stream_conv2d_25_source_start;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_802 <= _tmp_801;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_803 <= _tmp_802;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_804 <= _tmp_803;
      end 
      if(_stream_conv2d_25_stream_oready && _tmp_804) begin
        __variable_wdata_281 <= 0;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_807 <= _tmp_806;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_810 <= _tmp_809;
      end 
      if(_stream_conv2d_25_stream_oready && _tmp_810) begin
        __variable_wdata_281 <= 1;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_811 <= _stream_conv2d_25_source_start;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_812 <= _tmp_811;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_813 <= _tmp_812;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_814 <= _tmp_813;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_815 <= _tmp_814;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_816 <= _tmp_815;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_817 <= _tmp_816;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_818 <= _tmp_817;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_819 <= _tmp_818;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_820 <= _tmp_819;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_821 <= _tmp_820;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_822 <= _tmp_821;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_823 <= _tmp_822;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_824 <= _tmp_823;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_825 <= _tmp_824;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_826 <= _tmp_825;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_827 <= _tmp_826;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_828 <= _tmp_827;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_829 <= _tmp_828;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_830 <= _tmp_829;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_831 <= _tmp_830;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_832 <= _tmp_831;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_833 <= _tmp_832;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_834 <= _tmp_833;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_835 <= _tmp_834;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_836 <= _tmp_835;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_837 <= _tmp_836;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_838 <= _tmp_837;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_839 <= _tmp_838;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_840 <= _tmp_839;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_841 <= _tmp_840;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_842 <= _tmp_841;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_843 <= _tmp_842;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_844 <= _tmp_843;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_845 <= _tmp_844;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_846 <= _tmp_845;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_847 <= _stream_conv2d_25_source_stop;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_848 <= _tmp_847;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_849 <= _tmp_848;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_850 <= _tmp_849;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_851 <= _tmp_850;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_852 <= _tmp_851;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_853 <= _tmp_852;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_854 <= _tmp_853;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_855 <= _tmp_854;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_856 <= _tmp_855;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_857 <= _tmp_856;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_858 <= _tmp_857;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_859 <= _tmp_858;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_860 <= _tmp_859;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_861 <= _tmp_860;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_862 <= _tmp_861;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_863 <= _tmp_862;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_864 <= _tmp_863;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_865 <= _tmp_864;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_866 <= _tmp_865;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_867 <= _tmp_866;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_868 <= _tmp_867;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_869 <= _tmp_868;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_870 <= _tmp_869;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_871 <= _tmp_870;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_872 <= _tmp_871;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_873 <= _tmp_872;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_874 <= _tmp_873;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_875 <= _tmp_874;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_876 <= _tmp_875;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_877 <= _tmp_876;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_878 <= _tmp_877;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_879 <= _tmp_878;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_880 <= _tmp_879;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_881 <= _tmp_880;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_882 <= _tmp_881;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_883 <= _stream_conv2d_25_source_busy;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_884 <= _tmp_883;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_885 <= _tmp_884;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_886 <= _tmp_885;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_887 <= _tmp_886;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_888 <= _tmp_887;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_889 <= _tmp_888;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_890 <= _tmp_889;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_891 <= _tmp_890;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_892 <= _tmp_891;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_893 <= _tmp_892;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_894 <= _tmp_893;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_895 <= _tmp_894;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_896 <= _tmp_895;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_897 <= _tmp_896;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_898 <= _tmp_897;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_899 <= _tmp_898;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_900 <= _tmp_899;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_901 <= _tmp_900;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_902 <= _tmp_901;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_903 <= _tmp_902;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_904 <= _tmp_903;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_905 <= _tmp_904;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_906 <= _tmp_905;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_907 <= _tmp_906;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_908 <= _tmp_907;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_909 <= _tmp_908;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_910 <= _tmp_909;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_911 <= _tmp_910;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_912 <= _tmp_911;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_913 <= _tmp_912;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_914 <= _tmp_913;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_915 <= _tmp_914;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_916 <= _tmp_915;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_917 <= _tmp_916;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_918 <= _tmp_917;
      end 
      if(_stream_conv2d_25_stream_oready) begin
        _tmp_919 <= _stream_conv2d_25_sink_busy;
      end 
      if(!_stream_conv2d_25_sink_busy && _tmp_919) begin
        _stream_conv2d_25_busy_reg <= 0;
      end 
      if(_stream_conv2d_25_source_busy) begin
        _stream_conv2d_25_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_conv2d_25_fsm_1 = 1;
  localparam _stream_conv2d_25_fsm_2 = 2;
  localparam _stream_conv2d_25_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_fsm <= _stream_conv2d_25_fsm_init;
      _stream_conv2d_25_source_start <= 0;
      _stream_conv2d_25_source_busy <= 0;
      _stream_conv2d_25_stream_ivalid <= 0;
    end else begin
      if(_stream_conv2d_25_stream_oready && _tmp_797) begin
        _stream_conv2d_25_stream_ivalid <= 1;
      end 
      if(_stream_conv2d_25_stream_oready && _tmp_807) begin
        _stream_conv2d_25_stream_ivalid <= 0;
      end 
      case(_stream_conv2d_25_fsm)
        _stream_conv2d_25_fsm_init: begin
          if(_stream_conv2d_25_run_flag) begin
            _stream_conv2d_25_source_start <= 1;
          end 
          if(_stream_conv2d_25_run_flag) begin
            _stream_conv2d_25_fsm <= _stream_conv2d_25_fsm_1;
          end 
        end
        _stream_conv2d_25_fsm_1: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_start <= 0;
            _stream_conv2d_25_source_busy <= 1;
          end 
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_fsm <= _stream_conv2d_25_fsm_2;
          end 
        end
        _stream_conv2d_25_fsm_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_fsm <= _stream_conv2d_25_fsm_3;
          end 
        end
        _stream_conv2d_25_fsm_3: begin
          if(_stream_conv2d_25_stream_oready && (_stream_conv2d_25_source_11_idle && _stream_conv2d_25_source_13_idle && _stream_conv2d_25_source_15_idle && _stream_conv2d_25_source_20_idle && _stream_conv2d_25_source_21_idle && _stream_conv2d_25_source_22_idle && _stream_conv2d_25_source_23_idle && _stream_conv2d_25_source_24_idle && _stream_conv2d_25_source_25_idle && _stream_conv2d_25_source_26_idle && _stream_conv2d_25_source_27_idle && _stream_conv2d_25_source_28_idle && _stream_conv2d_25_source_29_idle && _stream_conv2d_25_source_30_idle && _stream_conv2d_25_source_31_idle && _stream_conv2d_25_source_32_idle && _stream_conv2d_25_source_33_idle && _stream_conv2d_25_source_34_idle && _stream_conv2d_25_source_35_idle && _stream_conv2d_25_source_36_idle && _stream_conv2d_25_source_37_idle && _stream_conv2d_25_source_7_idle && _stream_conv2d_25_source_9_idle && (_stream_conv2d_25_fsm == 3))) begin
            _stream_conv2d_25_source_busy <= 0;
          end 
          if(_stream_conv2d_25_stream_oready && (_stream_conv2d_25_source_11_idle && _stream_conv2d_25_source_13_idle && _stream_conv2d_25_source_15_idle && _stream_conv2d_25_source_20_idle && _stream_conv2d_25_source_21_idle && _stream_conv2d_25_source_22_idle && _stream_conv2d_25_source_23_idle && _stream_conv2d_25_source_24_idle && _stream_conv2d_25_source_25_idle && _stream_conv2d_25_source_26_idle && _stream_conv2d_25_source_27_idle && _stream_conv2d_25_source_28_idle && _stream_conv2d_25_source_29_idle && _stream_conv2d_25_source_30_idle && _stream_conv2d_25_source_31_idle && _stream_conv2d_25_source_32_idle && _stream_conv2d_25_source_33_idle && _stream_conv2d_25_source_34_idle && _stream_conv2d_25_source_35_idle && _stream_conv2d_25_source_36_idle && _stream_conv2d_25_source_37_idle && _stream_conv2d_25_source_7_idle && _stream_conv2d_25_source_9_idle && (_stream_conv2d_25_fsm == 3)) && _stream_conv2d_25_run_flag) begin
            _stream_conv2d_25_source_start <= 1;
          end 
          if(_stream_conv2d_25_stream_oready && (_stream_conv2d_25_source_11_idle && _stream_conv2d_25_source_13_idle && _stream_conv2d_25_source_15_idle && _stream_conv2d_25_source_20_idle && _stream_conv2d_25_source_21_idle && _stream_conv2d_25_source_22_idle && _stream_conv2d_25_source_23_idle && _stream_conv2d_25_source_24_idle && _stream_conv2d_25_source_25_idle && _stream_conv2d_25_source_26_idle && _stream_conv2d_25_source_27_idle && _stream_conv2d_25_source_28_idle && _stream_conv2d_25_source_29_idle && _stream_conv2d_25_source_30_idle && _stream_conv2d_25_source_31_idle && _stream_conv2d_25_source_32_idle && _stream_conv2d_25_source_33_idle && _stream_conv2d_25_source_34_idle && _stream_conv2d_25_source_35_idle && _stream_conv2d_25_source_36_idle && _stream_conv2d_25_source_37_idle && _stream_conv2d_25_source_7_idle && _stream_conv2d_25_source_9_idle && (_stream_conv2d_25_fsm == 3))) begin
            _stream_conv2d_25_fsm <= _stream_conv2d_25_fsm_init;
          end 
          if(_stream_conv2d_25_stream_oready && (_stream_conv2d_25_source_11_idle && _stream_conv2d_25_source_13_idle && _stream_conv2d_25_source_15_idle && _stream_conv2d_25_source_20_idle && _stream_conv2d_25_source_21_idle && _stream_conv2d_25_source_22_idle && _stream_conv2d_25_source_23_idle && _stream_conv2d_25_source_24_idle && _stream_conv2d_25_source_25_idle && _stream_conv2d_25_source_26_idle && _stream_conv2d_25_source_27_idle && _stream_conv2d_25_source_28_idle && _stream_conv2d_25_source_29_idle && _stream_conv2d_25_source_30_idle && _stream_conv2d_25_source_31_idle && _stream_conv2d_25_source_32_idle && _stream_conv2d_25_source_33_idle && _stream_conv2d_25_source_34_idle && _stream_conv2d_25_source_35_idle && _stream_conv2d_25_source_36_idle && _stream_conv2d_25_source_37_idle && _stream_conv2d_25_source_7_idle && _stream_conv2d_25_source_9_idle && (_stream_conv2d_25_fsm == 3)) && _stream_conv2d_25_run_flag) begin
            _stream_conv2d_25_fsm <= _stream_conv2d_25_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_27_source_1_source_ram_renable <= 0;
      _stream_max_pool_serial_27_source_1_source_fifo_deq <= 0;
      _stream_max_pool_serial_27_source_1_idle <= 1;
      _stream_max_pool_serial_27_sink_5_sink_wenable <= 0;
      _stream_max_pool_serial_27_sink_5_sink_fifo_enq <= 0;
      _stream_max_pool_serial_27_sink_6_sink_wenable <= 0;
      _stream_max_pool_serial_27_sink_6_sink_fifo_enq <= 0;
      __stream_max_pool_serial_27_stream_ivalid_1 <= 0;
      __stream_max_pool_serial_27_stream_ivalid_2 <= 0;
      __stream_max_pool_serial_27_stream_ivalid_3 <= 0;
      __stream_max_pool_serial_27_stream_ivalid_4 <= 0;
      __stream_max_pool_serial_27_stream_ivalid_5 <= 0;
      _counter_data_884 <= 1'sd0;
      _counter_count_884 <= 1'sd0;
      __delay_data_1123__variable_882 <= 0;
      __delay_data_1124_reinterpretcast_892 <= 0;
      __delay_data_1126__variable_883 <= 0;
      __delay_data_1129__variable_880 <= 0;
      _pointer_data_887 <= 0;
      __delay_data_1125__delay_1124_reinterpretcast_892 <= 0;
      __delay_data_1127__delay_1126__variable_883 <= 0;
      __delay_data_1130__delay_1129__variable_880 <= 0;
      _cond_data_894 <= 0;
      __delay_data_1128__delay_1127__delay_1126__variable_883 <= 0;
      __delay_data_1131__delay_1130__delay_1129__variable_880 <= 0;
      _stream_max_pool_serial_27_parameter_0_next_parameter_data <= 0;
      __variable_wdata_880 <= 0;
      _stream_max_pool_serial_27_parameter_2_next_parameter_data <= 0;
      __variable_wdata_882 <= 0;
      _stream_max_pool_serial_27_source_1_source_mode <= 5'b0;
      _stream_max_pool_serial_27_source_1_source_offset <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_size_0 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_stride_0 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_size_1 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_stride_1 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_size_2 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_stride_2 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_size_3 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_stride_3 <= 0;
      _stream_max_pool_serial_27_source_1_source_sel <= 0;
      _stream_max_pool_serial_27_source_1_source_offset_buf <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_cur_offset_0 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_cur_offset_1 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_cur_offset_2 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_cur_offset_3 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_count_0 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_count_1 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_count_2 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_count_3 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_size_buf_0 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_size_buf_1 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_size_buf_2 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_size_buf_3 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_stride_buf_0 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_stride_buf_1 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_stride_buf_2 <= 0;
      _source_stream_max_pool_serial_27_source_1_pat_stride_buf_3 <= 0;
      __variable_wdata_881 <= 0;
      _stream_max_pool_serial_27_source_1_source_ram_raddr <= 0;
      _tmp_972 <= 0;
      _tmp_973 <= 0;
      _tmp_974 <= 0;
      _tmp_975 <= 0;
      _tmp_976 <= 0;
      _tmp_977 <= 0;
      _tmp_978 <= 0;
      _tmp_981 <= 0;
      _tmp_982 <= 0;
      _tmp_983 <= 0;
      _tmp_984 <= 0;
      _tmp_985 <= 0;
      _tmp_986 <= 0;
      _tmp_987 <= 0;
      _tmp_988 <= 0;
      _tmp_989 <= 0;
      _tmp_990 <= 0;
      _tmp_991 <= 0;
      _tmp_992 <= 0;
      _tmp_993 <= 0;
      _tmp_994 <= 0;
      _stream_max_pool_serial_27_sink_5_sink_mode <= 5'b0;
      _stream_max_pool_serial_27_sink_5_sink_offset <= 0;
      _stream_max_pool_serial_27_sink_5_sink_size <= 0;
      _stream_max_pool_serial_27_sink_5_sink_stride <= 0;
      _stream_max_pool_serial_27_sink_5_sink_sel <= 0;
      _stream_max_pool_serial_27_sink_5_sink_offset_buf <= 0;
      _stream_max_pool_serial_27_sink_5_sink_size_buf <= 0;
      _stream_max_pool_serial_27_sink_5_sink_stride_buf <= 0;
      _stream_max_pool_serial_27_sink_5_sink_waddr <= 0;
      _stream_max_pool_serial_27_sink_5_sink_count <= 0;
      _stream_max_pool_serial_27_sink_5_sink_wdata <= 0;
      _tmp_1016 <= 0;
      _tmp_1017 <= 0;
      _tmp_1018 <= 0;
      _tmp_1019 <= 0;
      _tmp_1020 <= 0;
      _tmp_1021 <= 0;
      __variable_wdata_883 <= 0;
      _tmp_1022 <= 0;
      _tmp_1023 <= 0;
      _tmp_1024 <= 0;
      _tmp_1025 <= 0;
      _tmp_1028 <= 0;
      _tmp_1031 <= 0;
      _tmp_1032 <= 0;
      _tmp_1033 <= 0;
      _tmp_1034 <= 0;
      _tmp_1035 <= 0;
      _tmp_1036 <= 0;
      _tmp_1037 <= 0;
      _tmp_1038 <= 0;
      _tmp_1039 <= 0;
      _tmp_1040 <= 0;
      _tmp_1041 <= 0;
      _tmp_1042 <= 0;
      _tmp_1043 <= 0;
      _tmp_1044 <= 0;
      _tmp_1045 <= 0;
      _tmp_1046 <= 0;
      _tmp_1047 <= 0;
      _tmp_1048 <= 0;
      _tmp_1049 <= 0;
      _tmp_1050 <= 0;
      _tmp_1051 <= 0;
      _tmp_1052 <= 0;
      _tmp_1053 <= 0;
      _stream_max_pool_serial_27_busy_reg <= 0;
    end else begin
      if(_stream_max_pool_serial_27_stream_oready) begin
        _stream_max_pool_serial_27_source_1_source_ram_renable <= 0;
        _stream_max_pool_serial_27_source_1_source_fifo_deq <= 0;
      end 
      _stream_max_pool_serial_27_source_1_idle <= _stream_max_pool_serial_27_source_1_idle;
      if(_stream_max_pool_serial_27_stream_oready) begin
        _stream_max_pool_serial_27_sink_5_sink_wenable <= 0;
        _stream_max_pool_serial_27_sink_5_sink_fifo_enq <= 0;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _stream_max_pool_serial_27_sink_6_sink_wenable <= 0;
        _stream_max_pool_serial_27_sink_6_sink_fifo_enq <= 0;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        __stream_max_pool_serial_27_stream_ivalid_1 <= _stream_max_pool_serial_27_stream_ivalid;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        __stream_max_pool_serial_27_stream_ivalid_2 <= __stream_max_pool_serial_27_stream_ivalid_1;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        __stream_max_pool_serial_27_stream_ivalid_3 <= __stream_max_pool_serial_27_stream_ivalid_2;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        __stream_max_pool_serial_27_stream_ivalid_4 <= __stream_max_pool_serial_27_stream_ivalid_3;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        __stream_max_pool_serial_27_stream_ivalid_5 <= __stream_max_pool_serial_27_stream_ivalid_4;
      end 
      if(_stream_max_pool_serial_27_stream_ivalid && _stream_max_pool_serial_27_stream_oready && _counter_reset_cond_884) begin
        _counter_data_884 <= 1'sd0;
      end 
      if(_stream_max_pool_serial_27_stream_ivalid && _stream_max_pool_serial_27_stream_oready) begin
        _counter_data_884 <= _counter_current_count_884;
      end 
      if(_stream_max_pool_serial_27_stream_ivalid && _stream_max_pool_serial_27_stream_oready) begin
        _counter_count_884 <= (_counter_current_count_884 >= stream_max_pool_serial_27_parameter_0_data - 2'sd1)? _counter_current_count_884 + 2'sd1 - stream_max_pool_serial_27_parameter_0_data : _counter_current_count_884 + 2'sd1;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        __delay_data_1123__variable_882 <= stream_max_pool_serial_27_parameter_2_data;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        __delay_data_1124_reinterpretcast_892 <= _reinterpretcast_data_892;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        __delay_data_1126__variable_883 <= stream_max_pool_serial_27__reduce_reset_data;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        __delay_data_1129__variable_880 <= stream_max_pool_serial_27_parameter_0_data;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _pointer_data_887 <= __delay_data_1123__variable_882[_counter_data_884];
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        __delay_data_1125__delay_1124_reinterpretcast_892 <= __delay_data_1124_reinterpretcast_892;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        __delay_data_1127__delay_1126__variable_883 <= __delay_data_1126__variable_883;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        __delay_data_1130__delay_1129__variable_880 <= __delay_data_1129__variable_880;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _cond_data_894 <= (_pointer_data_887)? -33'sd2147483648 : __delay_data_1125__delay_1124_reinterpretcast_892;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        __delay_data_1128__delay_1127__delay_1126__variable_883 <= __delay_data_1127__delay_1126__variable_883;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        __delay_data_1131__delay_1130__delay_1129__variable_880 <= __delay_data_1130__delay_1129__variable_880;
      end 
      if(_set_flag_966) begin
        _stream_max_pool_serial_27_parameter_0_next_parameter_data <= 4;
      end 
      if(_stream_max_pool_serial_27_source_start) begin
        __variable_wdata_880 <= _stream_max_pool_serial_27_parameter_0_next_parameter_data;
      end 
      if(_set_flag_967) begin
        _stream_max_pool_serial_27_parameter_2_next_parameter_data <= max_pool_serial_27_stream_pad_masks;
      end 
      if(_stream_max_pool_serial_27_source_start) begin
        __variable_wdata_882 <= _stream_max_pool_serial_27_parameter_2_next_parameter_data;
      end 
      if(_set_flag_968) begin
        _stream_max_pool_serial_27_source_1_source_mode <= 5'b10;
        _stream_max_pool_serial_27_source_1_source_offset <= max_pool_serial_27_stream_act_local + max_pool_serial_27_act_page_comp_offset_buf;
      end 
      if(_set_flag_968) begin
        _source_stream_max_pool_serial_27_source_1_pat_size_0 <= 2;
        _source_stream_max_pool_serial_27_source_1_pat_stride_0 <= cparam_max_pool_serial_27_act_read_block;
      end 
      if(_set_flag_968) begin
        _source_stream_max_pool_serial_27_source_1_pat_size_1 <= 2;
        _source_stream_max_pool_serial_27_source_1_pat_stride_1 <= cparam_max_pool_serial_27_act_read_size;
      end 
      if(_set_flag_968) begin
        _source_stream_max_pool_serial_27_source_1_pat_size_2 <= cparam_max_pool_serial_27_stream_size;
        _source_stream_max_pool_serial_27_source_1_pat_stride_2 <= 1;
      end 
      if(_set_flag_968) begin
        _source_stream_max_pool_serial_27_source_1_pat_size_3 <= 1;
        _source_stream_max_pool_serial_27_source_1_pat_stride_3 <= 0;
      end 
      if(_set_flag_968) begin
        _stream_max_pool_serial_27_source_1_source_sel <= 1;
      end 
      if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
        _stream_max_pool_serial_27_source_1_source_offset_buf <= _stream_max_pool_serial_27_source_1_source_offset;
      end 
      if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_cur_offset_0 <= 0;
      end 
      if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_cur_offset_1 <= 0;
      end 
      if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_cur_offset_2 <= 0;
      end 
      if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_cur_offset_3 <= 0;
      end 
      if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_count_0 <= _source_stream_max_pool_serial_27_source_1_pat_size_0 - 1;
      end 
      if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_count_1 <= _source_stream_max_pool_serial_27_source_1_pat_size_1 - 1;
      end 
      if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_count_2 <= _source_stream_max_pool_serial_27_source_1_pat_size_2 - 1;
      end 
      if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_count_3 <= _source_stream_max_pool_serial_27_source_1_pat_size_3 - 1;
      end 
      if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_size_buf_0 <= _source_stream_max_pool_serial_27_source_1_pat_size_0;
      end 
      if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_size_buf_1 <= _source_stream_max_pool_serial_27_source_1_pat_size_1;
      end 
      if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_size_buf_2 <= _source_stream_max_pool_serial_27_source_1_pat_size_2;
      end 
      if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_size_buf_3 <= _source_stream_max_pool_serial_27_source_1_pat_size_3;
      end 
      if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_stride_buf_0 <= _source_stream_max_pool_serial_27_source_1_pat_stride_0;
      end 
      if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_stride_buf_1 <= _source_stream_max_pool_serial_27_source_1_pat_stride_1;
      end 
      if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_stride_buf_2 <= _source_stream_max_pool_serial_27_source_1_pat_stride_2;
      end 
      if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_stride_buf_3 <= _source_stream_max_pool_serial_27_source_1_pat_stride_3;
      end 
      if(_stream_max_pool_serial_27_stream_oready && _stream_max_pool_serial_27_source_busy && _stream_max_pool_serial_27_is_root) begin
        __variable_wdata_881 <= _stream_max_pool_serial_27_source_1_source_ram_rdata;
      end 
      if((_stream_max_pool_serial_27_source_1_source_pat_fsm_0 == 1) && _stream_max_pool_serial_27_stream_oready) begin
        _stream_max_pool_serial_27_source_1_idle <= 0;
        _stream_max_pool_serial_27_source_1_source_ram_raddr <= _stream_max_pool_serial_27_source_1_source_pat_all_offset;
        _stream_max_pool_serial_27_source_1_source_ram_renable <= 1;
      end 
      if((_stream_max_pool_serial_27_source_1_source_pat_fsm_0 == 1) && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_cur_offset_0 <= _source_stream_max_pool_serial_27_source_1_pat_cur_offset_0 + _source_stream_max_pool_serial_27_source_1_pat_stride_buf_0;
        _source_stream_max_pool_serial_27_source_1_pat_count_0 <= _source_stream_max_pool_serial_27_source_1_pat_count_0 - 1;
      end 
      if((_stream_max_pool_serial_27_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_27_source_1_pat_count_0 == 0) && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_cur_offset_0 <= 0;
        _source_stream_max_pool_serial_27_source_1_pat_count_0 <= _source_stream_max_pool_serial_27_source_1_pat_size_buf_0 - 1;
      end 
      if((_stream_max_pool_serial_27_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_27_source_1_pat_count_0 == 0) && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_cur_offset_1 <= _source_stream_max_pool_serial_27_source_1_pat_cur_offset_1 + _source_stream_max_pool_serial_27_source_1_pat_stride_buf_1;
        _source_stream_max_pool_serial_27_source_1_pat_count_1 <= _source_stream_max_pool_serial_27_source_1_pat_count_1 - 1;
      end 
      if((_stream_max_pool_serial_27_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_27_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_27_source_1_pat_count_1 == 0) && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_cur_offset_1 <= 0;
        _source_stream_max_pool_serial_27_source_1_pat_count_1 <= _source_stream_max_pool_serial_27_source_1_pat_size_buf_1 - 1;
      end 
      if((_stream_max_pool_serial_27_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_27_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_27_source_1_pat_count_1 == 0)) && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_cur_offset_2 <= _source_stream_max_pool_serial_27_source_1_pat_cur_offset_2 + _source_stream_max_pool_serial_27_source_1_pat_stride_buf_2;
        _source_stream_max_pool_serial_27_source_1_pat_count_2 <= _source_stream_max_pool_serial_27_source_1_pat_count_2 - 1;
      end 
      if((_stream_max_pool_serial_27_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_27_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_27_source_1_pat_count_1 == 0)) && (_source_stream_max_pool_serial_27_source_1_pat_count_2 == 0) && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_cur_offset_2 <= 0;
        _source_stream_max_pool_serial_27_source_1_pat_count_2 <= _source_stream_max_pool_serial_27_source_1_pat_size_buf_2 - 1;
      end 
      if((_stream_max_pool_serial_27_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_27_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_27_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_27_source_1_pat_count_2 == 0)) && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_cur_offset_3 <= _source_stream_max_pool_serial_27_source_1_pat_cur_offset_3 + _source_stream_max_pool_serial_27_source_1_pat_stride_buf_3;
        _source_stream_max_pool_serial_27_source_1_pat_count_3 <= _source_stream_max_pool_serial_27_source_1_pat_count_3 - 1;
      end 
      if((_stream_max_pool_serial_27_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_27_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_27_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_27_source_1_pat_count_2 == 0)) && (_source_stream_max_pool_serial_27_source_1_pat_count_3 == 0) && _stream_max_pool_serial_27_stream_oready) begin
        _source_stream_max_pool_serial_27_source_1_pat_cur_offset_3 <= 0;
        _source_stream_max_pool_serial_27_source_1_pat_count_3 <= _source_stream_max_pool_serial_27_source_1_pat_size_buf_3 - 1;
      end 
      if((_stream_max_pool_serial_27_source_1_source_pat_fsm_0 == 1) && _stream_max_pool_serial_27_source_stop && _stream_max_pool_serial_27_stream_oready) begin
        _stream_max_pool_serial_27_source_1_source_ram_renable <= 0;
        _stream_max_pool_serial_27_source_1_idle <= 1;
      end 
      if((_stream_max_pool_serial_27_source_1_source_pat_fsm_0 == 2) && _stream_max_pool_serial_27_stream_oready) begin
        _stream_max_pool_serial_27_source_1_source_ram_renable <= 0;
        _stream_max_pool_serial_27_source_1_idle <= 1;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_972 <= _set_flag_971;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_973 <= _tmp_972;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_974 <= _tmp_973;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_975 <= _tmp_974;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_976 <= _tmp_975;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_977 <= _tmp_976;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_978 <= _tmp_977;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_981 <= _tmp_980;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_982 <= _tmp_981;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_983 <= _tmp_982;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_984 <= _tmp_983;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_985 <= _tmp_984;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_986 <= _tmp_985;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_987 <= _tmp_986;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_988 <= cparam_max_pool_serial_27_stream_size;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_989 <= _tmp_988;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_990 <= _tmp_989;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_991 <= _tmp_990;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_992 <= _tmp_991;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_993 <= _tmp_992;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_994 <= _tmp_993;
      end 
      if(_tmp_978) begin
        _stream_max_pool_serial_27_sink_5_sink_mode <= 5'b1;
        _stream_max_pool_serial_27_sink_5_sink_offset <= _tmp_987;
        _stream_max_pool_serial_27_sink_5_sink_size <= _tmp_994;
        _stream_max_pool_serial_27_sink_5_sink_stride <= 1;
      end 
      if(_tmp_978) begin
        _stream_max_pool_serial_27_sink_5_sink_sel <= 2;
      end 
      if(_stream_max_pool_serial_27_sink_start && _stream_max_pool_serial_27_sink_5_sink_mode & 5'b1 && _stream_max_pool_serial_27_stream_oready) begin
        _stream_max_pool_serial_27_sink_5_sink_offset_buf <= _stream_max_pool_serial_27_sink_5_sink_offset;
        _stream_max_pool_serial_27_sink_5_sink_size_buf <= _stream_max_pool_serial_27_sink_5_sink_size;
        _stream_max_pool_serial_27_sink_5_sink_stride_buf <= _stream_max_pool_serial_27_sink_5_sink_stride;
      end 
      if((_stream_max_pool_serial_27_sink_5_sink_fsm_1 == 1) && _stream_max_pool_serial_27_stream_oready) begin
        _stream_max_pool_serial_27_sink_5_sink_waddr <= _stream_max_pool_serial_27_sink_5_sink_offset_buf - _stream_max_pool_serial_27_sink_5_sink_stride_buf;
        _stream_max_pool_serial_27_sink_5_sink_count <= _stream_max_pool_serial_27_sink_5_sink_size_buf;
      end 
      if((_stream_max_pool_serial_27_sink_5_sink_fsm_1 == 2) && stream_max_pool_serial_27_sink_6_data && _stream_max_pool_serial_27_stream_oready) begin
        _stream_max_pool_serial_27_sink_5_sink_waddr <= _stream_max_pool_serial_27_sink_5_sink_waddr + _stream_max_pool_serial_27_sink_5_sink_stride_buf;
        _stream_max_pool_serial_27_sink_5_sink_wdata <= stream_max_pool_serial_27_sink_5_data;
        _stream_max_pool_serial_27_sink_5_sink_wenable <= 1;
        _stream_max_pool_serial_27_sink_5_sink_count <= _stream_max_pool_serial_27_sink_5_sink_count - 1;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1016 <= _stream_max_pool_serial_27_source_start;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1017 <= _tmp_1016;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1018 <= _tmp_1017;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1019 <= _stream_max_pool_serial_27_source_start;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1020 <= _tmp_1019;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1021 <= _tmp_1020;
      end 
      if(_stream_max_pool_serial_27_stream_oready && _tmp_1021) begin
        __variable_wdata_883 <= 1;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1022 <= _stream_max_pool_serial_27_source_start;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1023 <= _tmp_1022;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1024 <= _tmp_1023;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1025 <= _tmp_1024;
      end 
      if(_stream_max_pool_serial_27_stream_oready && _tmp_1025) begin
        __variable_wdata_883 <= 0;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1028 <= _tmp_1027;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1031 <= _tmp_1030;
      end 
      if(_stream_max_pool_serial_27_stream_oready && _tmp_1031) begin
        __variable_wdata_883 <= 1;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1032 <= _stream_max_pool_serial_27_source_start;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1033 <= _tmp_1032;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1034 <= _tmp_1033;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1035 <= _tmp_1034;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1036 <= _tmp_1035;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1037 <= _tmp_1036;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1038 <= _tmp_1037;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1039 <= _stream_max_pool_serial_27_source_stop;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1040 <= _tmp_1039;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1041 <= _tmp_1040;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1042 <= _tmp_1041;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1043 <= _tmp_1042;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1044 <= _tmp_1043;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1045 <= _tmp_1044;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1046 <= _stream_max_pool_serial_27_source_busy;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1047 <= _tmp_1046;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1048 <= _tmp_1047;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1049 <= _tmp_1048;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1050 <= _tmp_1049;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1051 <= _tmp_1050;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1052 <= _tmp_1051;
      end 
      if(_stream_max_pool_serial_27_stream_oready) begin
        _tmp_1053 <= _stream_max_pool_serial_27_sink_busy;
      end 
      if(!_stream_max_pool_serial_27_sink_busy && _tmp_1053) begin
        _stream_max_pool_serial_27_busy_reg <= 0;
      end 
      if(_stream_max_pool_serial_27_source_busy) begin
        _stream_max_pool_serial_27_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_max_pool_serial_27_fsm_1 = 1;
  localparam _stream_max_pool_serial_27_fsm_2 = 2;
  localparam _stream_max_pool_serial_27_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_27_fsm <= _stream_max_pool_serial_27_fsm_init;
      _stream_max_pool_serial_27_source_start <= 0;
      _stream_max_pool_serial_27_source_busy <= 0;
      _stream_max_pool_serial_27_stream_ivalid <= 0;
    end else begin
      if(_stream_max_pool_serial_27_stream_oready && _tmp_1018) begin
        _stream_max_pool_serial_27_stream_ivalid <= 1;
      end 
      if(_stream_max_pool_serial_27_stream_oready && _tmp_1028) begin
        _stream_max_pool_serial_27_stream_ivalid <= 0;
      end 
      case(_stream_max_pool_serial_27_fsm)
        _stream_max_pool_serial_27_fsm_init: begin
          if(_stream_max_pool_serial_27_run_flag) begin
            _stream_max_pool_serial_27_source_start <= 1;
          end 
          if(_stream_max_pool_serial_27_run_flag) begin
            _stream_max_pool_serial_27_fsm <= _stream_max_pool_serial_27_fsm_1;
          end 
        end
        _stream_max_pool_serial_27_fsm_1: begin
          if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_stream_oready) begin
            _stream_max_pool_serial_27_source_start <= 0;
            _stream_max_pool_serial_27_source_busy <= 1;
          end 
          if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_stream_oready) begin
            _stream_max_pool_serial_27_fsm <= _stream_max_pool_serial_27_fsm_2;
          end 
        end
        _stream_max_pool_serial_27_fsm_2: begin
          if(_stream_max_pool_serial_27_stream_oready) begin
            _stream_max_pool_serial_27_fsm <= _stream_max_pool_serial_27_fsm_3;
          end 
        end
        _stream_max_pool_serial_27_fsm_3: begin
          if(_stream_max_pool_serial_27_stream_oready && (_stream_max_pool_serial_27_source_1_idle && (_stream_max_pool_serial_27_fsm == 3))) begin
            _stream_max_pool_serial_27_source_busy <= 0;
          end 
          if(_stream_max_pool_serial_27_stream_oready && (_stream_max_pool_serial_27_source_1_idle && (_stream_max_pool_serial_27_fsm == 3)) && _stream_max_pool_serial_27_run_flag) begin
            _stream_max_pool_serial_27_source_start <= 1;
          end 
          if(_stream_max_pool_serial_27_stream_oready && (_stream_max_pool_serial_27_source_1_idle && (_stream_max_pool_serial_27_fsm == 3))) begin
            _stream_max_pool_serial_27_fsm <= _stream_max_pool_serial_27_fsm_init;
          end 
          if(_stream_max_pool_serial_27_stream_oready && (_stream_max_pool_serial_27_source_1_idle && (_stream_max_pool_serial_27_fsm == 3)) && _stream_max_pool_serial_27_run_flag) begin
            _stream_max_pool_serial_27_fsm <= _stream_max_pool_serial_27_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_47_source_1_source_ram_renable <= 0;
      _stream_max_pool_47_source_1_source_fifo_deq <= 0;
      _stream_max_pool_47_source_1_idle <= 1;
      _stream_max_pool_47_source_2_source_ram_renable <= 0;
      _stream_max_pool_47_source_2_source_fifo_deq <= 0;
      _stream_max_pool_47_source_2_idle <= 1;
      _stream_max_pool_47_source_3_source_ram_renable <= 0;
      _stream_max_pool_47_source_3_source_fifo_deq <= 0;
      _stream_max_pool_47_source_3_idle <= 1;
      _stream_max_pool_47_source_4_source_ram_renable <= 0;
      _stream_max_pool_47_source_4_source_fifo_deq <= 0;
      _stream_max_pool_47_source_4_idle <= 1;
      _stream_max_pool_47_sink_6_sink_wenable <= 0;
      _stream_max_pool_47_sink_6_sink_fifo_enq <= 0;
      __stream_max_pool_47_stream_ivalid_1 <= 0;
      __stream_max_pool_47_stream_ivalid_2 <= 0;
      __stream_max_pool_47_stream_ivalid_3 <= 0;
      __stream_max_pool_47_stream_ivalid_4 <= 0;
      __stream_max_pool_47_stream_ivalid_5 <= 0;
      __stream_max_pool_47_stream_ivalid_6 <= 0;
      _cond_data_927 <= 0;
      _cond_data_930 <= 0;
      _cond_data_933 <= 0;
      _cond_data_936 <= 0;
      _stream_max_pool_47_parameter_0_next_parameter_data <= 0;
      __variable_wdata_899 <= 0;
      _stream_max_pool_47_source_1_source_mode <= 5'b0;
      _stream_max_pool_47_source_1_source_offset <= 0;
      _stream_max_pool_47_source_1_source_size <= 0;
      _stream_max_pool_47_source_1_source_stride <= 0;
      _stream_max_pool_47_source_1_source_sel <= 0;
      _stream_max_pool_47_source_1_source_offset_buf <= 0;
      _stream_max_pool_47_source_1_source_size_buf <= 0;
      _stream_max_pool_47_source_1_source_stride_buf <= 0;
      __variable_wdata_900 <= 0;
      _stream_max_pool_47_source_1_source_ram_raddr <= 0;
      _stream_max_pool_47_source_1_source_count <= 0;
      _stream_max_pool_47_source_2_source_mode <= 5'b0;
      _stream_max_pool_47_source_2_source_offset <= 0;
      _stream_max_pool_47_source_2_source_size <= 0;
      _stream_max_pool_47_source_2_source_stride <= 0;
      _stream_max_pool_47_source_2_source_sel <= 0;
      _stream_max_pool_47_source_2_source_offset_buf <= 0;
      _stream_max_pool_47_source_2_source_size_buf <= 0;
      _stream_max_pool_47_source_2_source_stride_buf <= 0;
      __variable_wdata_901 <= 0;
      _stream_max_pool_47_source_2_source_ram_raddr <= 0;
      _stream_max_pool_47_source_2_source_count <= 0;
      _stream_max_pool_47_source_3_source_mode <= 5'b0;
      _stream_max_pool_47_source_3_source_offset <= 0;
      _stream_max_pool_47_source_3_source_size <= 0;
      _stream_max_pool_47_source_3_source_stride <= 0;
      _stream_max_pool_47_source_3_source_sel <= 0;
      _stream_max_pool_47_source_3_source_offset_buf <= 0;
      _stream_max_pool_47_source_3_source_size_buf <= 0;
      _stream_max_pool_47_source_3_source_stride_buf <= 0;
      __variable_wdata_902 <= 0;
      _stream_max_pool_47_source_3_source_ram_raddr <= 0;
      _stream_max_pool_47_source_3_source_count <= 0;
      _stream_max_pool_47_source_4_source_mode <= 5'b0;
      _stream_max_pool_47_source_4_source_offset <= 0;
      _stream_max_pool_47_source_4_source_size <= 0;
      _stream_max_pool_47_source_4_source_stride <= 0;
      _stream_max_pool_47_source_4_source_sel <= 0;
      _stream_max_pool_47_source_4_source_offset_buf <= 0;
      _stream_max_pool_47_source_4_source_size_buf <= 0;
      _stream_max_pool_47_source_4_source_stride_buf <= 0;
      __variable_wdata_903 <= 0;
      _stream_max_pool_47_source_4_source_ram_raddr <= 0;
      _stream_max_pool_47_source_4_source_count <= 0;
      _tmp_1114 <= 0;
      _tmp_1115 <= 0;
      _tmp_1116 <= 0;
      _tmp_1117 <= 0;
      _tmp_1118 <= 0;
      _tmp_1119 <= 0;
      _tmp_1120 <= 0;
      _tmp_1121 <= 0;
      _tmp_1124 <= 0;
      _tmp_1125 <= 0;
      _tmp_1126 <= 0;
      _tmp_1127 <= 0;
      _tmp_1128 <= 0;
      _tmp_1129 <= 0;
      _tmp_1130 <= 0;
      _tmp_1131 <= 0;
      _tmp_1132 <= 0;
      _tmp_1133 <= 0;
      _tmp_1134 <= 0;
      _tmp_1135 <= 0;
      _tmp_1136 <= 0;
      _tmp_1137 <= 0;
      _tmp_1138 <= 0;
      _tmp_1139 <= 0;
      _stream_max_pool_47_sink_6_sink_mode <= 5'b0;
      _stream_max_pool_47_sink_6_sink_offset <= 0;
      _stream_max_pool_47_sink_6_sink_size <= 0;
      _stream_max_pool_47_sink_6_sink_stride <= 0;
      _stream_max_pool_47_sink_6_sink_sel <= 0;
      _stream_max_pool_47_sink_6_sink_offset_buf <= 0;
      _stream_max_pool_47_sink_6_sink_size_buf <= 0;
      _stream_max_pool_47_sink_6_sink_stride_buf <= 0;
      _stream_max_pool_47_sink_6_sink_waddr <= 0;
      _stream_max_pool_47_sink_6_sink_count <= 0;
      _stream_max_pool_47_sink_6_sink_wdata <= 0;
      _tmp_1163 <= 0;
      _tmp_1164 <= 0;
      _tmp_1165 <= 0;
      _tmp_1168 <= 0;
      _tmp_1169 <= 0;
      _tmp_1170 <= 0;
      _tmp_1171 <= 0;
      _tmp_1172 <= 0;
      _tmp_1173 <= 0;
      _tmp_1174 <= 0;
      _tmp_1175 <= 0;
      _tmp_1176 <= 0;
      _tmp_1177 <= 0;
      _tmp_1178 <= 0;
      _tmp_1179 <= 0;
      _tmp_1180 <= 0;
      _tmp_1181 <= 0;
      _tmp_1182 <= 0;
      _tmp_1183 <= 0;
      _tmp_1184 <= 0;
      _tmp_1185 <= 0;
      _tmp_1186 <= 0;
      _tmp_1187 <= 0;
      _tmp_1188 <= 0;
      _tmp_1189 <= 0;
      _tmp_1190 <= 0;
      _tmp_1191 <= 0;
      _tmp_1192 <= 0;
      _tmp_1193 <= 0;
      _stream_max_pool_47_busy_reg <= 0;
    end else begin
      if(_stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_1_source_ram_renable <= 0;
        _stream_max_pool_47_source_1_source_fifo_deq <= 0;
      end 
      _stream_max_pool_47_source_1_idle <= _stream_max_pool_47_source_1_idle;
      if(_stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_2_source_ram_renable <= 0;
        _stream_max_pool_47_source_2_source_fifo_deq <= 0;
      end 
      _stream_max_pool_47_source_2_idle <= _stream_max_pool_47_source_2_idle;
      if(_stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_3_source_ram_renable <= 0;
        _stream_max_pool_47_source_3_source_fifo_deq <= 0;
      end 
      _stream_max_pool_47_source_3_idle <= _stream_max_pool_47_source_3_idle;
      if(_stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_4_source_ram_renable <= 0;
        _stream_max_pool_47_source_4_source_fifo_deq <= 0;
      end 
      _stream_max_pool_47_source_4_idle <= _stream_max_pool_47_source_4_idle;
      if(_stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_sink_6_sink_wenable <= 0;
        _stream_max_pool_47_sink_6_sink_fifo_enq <= 0;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        __stream_max_pool_47_stream_ivalid_1 <= _stream_max_pool_47_stream_ivalid;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        __stream_max_pool_47_stream_ivalid_2 <= __stream_max_pool_47_stream_ivalid_1;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        __stream_max_pool_47_stream_ivalid_3 <= __stream_max_pool_47_stream_ivalid_2;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        __stream_max_pool_47_stream_ivalid_4 <= __stream_max_pool_47_stream_ivalid_3;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        __stream_max_pool_47_stream_ivalid_5 <= __stream_max_pool_47_stream_ivalid_4;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        __stream_max_pool_47_stream_ivalid_6 <= __stream_max_pool_47_stream_ivalid_5;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _cond_data_927 <= (_pointer_data_925)? -33'sd2147483648 : _reinterpretcast_data_920;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _cond_data_930 <= (_pointer_data_928)? -33'sd2147483648 : _reinterpretcast_data_921;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _cond_data_933 <= (_pointer_data_931)? -33'sd2147483648 : _reinterpretcast_data_922;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _cond_data_936 <= (_pointer_data_934)? -33'sd2147483648 : _reinterpretcast_data_923;
      end 
      if(_set_flag_1100) begin
        _stream_max_pool_47_parameter_0_next_parameter_data <= max_pool_47_stream_pad_masks;
      end 
      if(_stream_max_pool_47_source_start) begin
        __variable_wdata_899 <= _stream_max_pool_47_parameter_0_next_parameter_data;
      end 
      if(_set_flag_1101) begin
        _stream_max_pool_47_source_1_source_mode <= 5'b1;
        _stream_max_pool_47_source_1_source_offset <= max_pool_47_stream_act_local_0 + max_pool_47_act_page_comp_offset_buf_0;
        _stream_max_pool_47_source_1_source_size <= cparam_max_pool_47_stream_size;
        _stream_max_pool_47_source_1_source_stride <= 1;
      end 
      if(_set_flag_1101) begin
        _stream_max_pool_47_source_1_source_sel <= 1;
      end 
      if(_stream_max_pool_47_source_start && _stream_max_pool_47_source_1_source_mode & 5'b1 && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_1_source_offset_buf <= _stream_max_pool_47_source_1_source_offset;
        _stream_max_pool_47_source_1_source_size_buf <= _stream_max_pool_47_source_1_source_size;
        _stream_max_pool_47_source_1_source_stride_buf <= _stream_max_pool_47_source_1_source_stride;
      end 
      if(_stream_max_pool_47_stream_oready && _stream_max_pool_47_source_busy && _stream_max_pool_47_is_root) begin
        __variable_wdata_900 <= _stream_max_pool_47_source_1_source_ram_rdata;
      end 
      if((_stream_max_pool_47_source_1_source_fsm_0 == 1) && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_1_idle <= 0;
        _stream_max_pool_47_source_1_source_ram_raddr <= _stream_max_pool_47_source_1_source_offset_buf;
        _stream_max_pool_47_source_1_source_ram_renable <= 1;
        _stream_max_pool_47_source_1_source_count <= _stream_max_pool_47_source_1_source_size_buf;
      end 
      if((_stream_max_pool_47_source_1_source_fsm_0 == 2) && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_1_source_ram_raddr <= _stream_max_pool_47_source_1_source_ram_raddr + _stream_max_pool_47_source_1_source_stride_buf;
        _stream_max_pool_47_source_1_source_ram_renable <= 1;
        _stream_max_pool_47_source_1_source_count <= _stream_max_pool_47_source_1_source_count - 1;
      end 
      if((_stream_max_pool_47_source_1_source_fsm_0 == 2) && (_stream_max_pool_47_source_1_source_count == 1) && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_1_source_ram_renable <= 0;
        _stream_max_pool_47_source_1_idle <= 1;
      end 
      if((_stream_max_pool_47_source_1_source_fsm_0 == 2) && _stream_max_pool_47_source_stop && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_1_source_ram_renable <= 0;
        _stream_max_pool_47_source_1_idle <= 1;
      end 
      if(_set_flag_1104) begin
        _stream_max_pool_47_source_2_source_mode <= 5'b1;
        _stream_max_pool_47_source_2_source_offset <= max_pool_47_stream_act_local_1 + max_pool_47_act_page_comp_offset_buf_0;
        _stream_max_pool_47_source_2_source_size <= cparam_max_pool_47_stream_size;
        _stream_max_pool_47_source_2_source_stride <= 1;
      end 
      if(_set_flag_1104) begin
        _stream_max_pool_47_source_2_source_sel <= 2;
      end 
      if(_stream_max_pool_47_source_start && _stream_max_pool_47_source_2_source_mode & 5'b1 && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_2_source_offset_buf <= _stream_max_pool_47_source_2_source_offset;
        _stream_max_pool_47_source_2_source_size_buf <= _stream_max_pool_47_source_2_source_size;
        _stream_max_pool_47_source_2_source_stride_buf <= _stream_max_pool_47_source_2_source_stride;
      end 
      if(_stream_max_pool_47_stream_oready && _stream_max_pool_47_source_busy && _stream_max_pool_47_is_root) begin
        __variable_wdata_901 <= _stream_max_pool_47_source_2_source_ram_rdata;
      end 
      if((_stream_max_pool_47_source_2_source_fsm_1 == 1) && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_2_idle <= 0;
        _stream_max_pool_47_source_2_source_ram_raddr <= _stream_max_pool_47_source_2_source_offset_buf;
        _stream_max_pool_47_source_2_source_ram_renable <= 1;
        _stream_max_pool_47_source_2_source_count <= _stream_max_pool_47_source_2_source_size_buf;
      end 
      if((_stream_max_pool_47_source_2_source_fsm_1 == 2) && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_2_source_ram_raddr <= _stream_max_pool_47_source_2_source_ram_raddr + _stream_max_pool_47_source_2_source_stride_buf;
        _stream_max_pool_47_source_2_source_ram_renable <= 1;
        _stream_max_pool_47_source_2_source_count <= _stream_max_pool_47_source_2_source_count - 1;
      end 
      if((_stream_max_pool_47_source_2_source_fsm_1 == 2) && (_stream_max_pool_47_source_2_source_count == 1) && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_2_source_ram_renable <= 0;
        _stream_max_pool_47_source_2_idle <= 1;
      end 
      if((_stream_max_pool_47_source_2_source_fsm_1 == 2) && _stream_max_pool_47_source_stop && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_2_source_ram_renable <= 0;
        _stream_max_pool_47_source_2_idle <= 1;
      end 
      if(_set_flag_1107) begin
        _stream_max_pool_47_source_3_source_mode <= 5'b1;
        _stream_max_pool_47_source_3_source_offset <= max_pool_47_stream_act_local_2 + max_pool_47_act_page_comp_offset_buf_1;
        _stream_max_pool_47_source_3_source_size <= cparam_max_pool_47_stream_size;
        _stream_max_pool_47_source_3_source_stride <= 1;
      end 
      if(_set_flag_1107) begin
        _stream_max_pool_47_source_3_source_sel <= 3;
      end 
      if(_stream_max_pool_47_source_start && _stream_max_pool_47_source_3_source_mode & 5'b1 && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_3_source_offset_buf <= _stream_max_pool_47_source_3_source_offset;
        _stream_max_pool_47_source_3_source_size_buf <= _stream_max_pool_47_source_3_source_size;
        _stream_max_pool_47_source_3_source_stride_buf <= _stream_max_pool_47_source_3_source_stride;
      end 
      if(_stream_max_pool_47_stream_oready && _stream_max_pool_47_source_busy && _stream_max_pool_47_is_root) begin
        __variable_wdata_902 <= _stream_max_pool_47_source_3_source_ram_rdata;
      end 
      if((_stream_max_pool_47_source_3_source_fsm_2 == 1) && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_3_idle <= 0;
        _stream_max_pool_47_source_3_source_ram_raddr <= _stream_max_pool_47_source_3_source_offset_buf;
        _stream_max_pool_47_source_3_source_ram_renable <= 1;
        _stream_max_pool_47_source_3_source_count <= _stream_max_pool_47_source_3_source_size_buf;
      end 
      if((_stream_max_pool_47_source_3_source_fsm_2 == 2) && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_3_source_ram_raddr <= _stream_max_pool_47_source_3_source_ram_raddr + _stream_max_pool_47_source_3_source_stride_buf;
        _stream_max_pool_47_source_3_source_ram_renable <= 1;
        _stream_max_pool_47_source_3_source_count <= _stream_max_pool_47_source_3_source_count - 1;
      end 
      if((_stream_max_pool_47_source_3_source_fsm_2 == 2) && (_stream_max_pool_47_source_3_source_count == 1) && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_3_source_ram_renable <= 0;
        _stream_max_pool_47_source_3_idle <= 1;
      end 
      if((_stream_max_pool_47_source_3_source_fsm_2 == 2) && _stream_max_pool_47_source_stop && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_3_source_ram_renable <= 0;
        _stream_max_pool_47_source_3_idle <= 1;
      end 
      if(_set_flag_1110) begin
        _stream_max_pool_47_source_4_source_mode <= 5'b1;
        _stream_max_pool_47_source_4_source_offset <= max_pool_47_stream_act_local_3 + max_pool_47_act_page_comp_offset_buf_1;
        _stream_max_pool_47_source_4_source_size <= cparam_max_pool_47_stream_size;
        _stream_max_pool_47_source_4_source_stride <= 1;
      end 
      if(_set_flag_1110) begin
        _stream_max_pool_47_source_4_source_sel <= 4;
      end 
      if(_stream_max_pool_47_source_start && _stream_max_pool_47_source_4_source_mode & 5'b1 && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_4_source_offset_buf <= _stream_max_pool_47_source_4_source_offset;
        _stream_max_pool_47_source_4_source_size_buf <= _stream_max_pool_47_source_4_source_size;
        _stream_max_pool_47_source_4_source_stride_buf <= _stream_max_pool_47_source_4_source_stride;
      end 
      if(_stream_max_pool_47_stream_oready && _stream_max_pool_47_source_busy && _stream_max_pool_47_is_root) begin
        __variable_wdata_903 <= _stream_max_pool_47_source_4_source_ram_rdata;
      end 
      if((_stream_max_pool_47_source_4_source_fsm_3 == 1) && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_4_idle <= 0;
        _stream_max_pool_47_source_4_source_ram_raddr <= _stream_max_pool_47_source_4_source_offset_buf;
        _stream_max_pool_47_source_4_source_ram_renable <= 1;
        _stream_max_pool_47_source_4_source_count <= _stream_max_pool_47_source_4_source_size_buf;
      end 
      if((_stream_max_pool_47_source_4_source_fsm_3 == 2) && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_4_source_ram_raddr <= _stream_max_pool_47_source_4_source_ram_raddr + _stream_max_pool_47_source_4_source_stride_buf;
        _stream_max_pool_47_source_4_source_ram_renable <= 1;
        _stream_max_pool_47_source_4_source_count <= _stream_max_pool_47_source_4_source_count - 1;
      end 
      if((_stream_max_pool_47_source_4_source_fsm_3 == 2) && (_stream_max_pool_47_source_4_source_count == 1) && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_4_source_ram_renable <= 0;
        _stream_max_pool_47_source_4_idle <= 1;
      end 
      if((_stream_max_pool_47_source_4_source_fsm_3 == 2) && _stream_max_pool_47_source_stop && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_source_4_source_ram_renable <= 0;
        _stream_max_pool_47_source_4_idle <= 1;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1114 <= _set_flag_1113;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1115 <= _tmp_1114;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1116 <= _tmp_1115;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1117 <= _tmp_1116;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1118 <= _tmp_1117;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1119 <= _tmp_1118;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1120 <= _tmp_1119;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1121 <= _tmp_1120;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1124 <= _tmp_1123;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1125 <= _tmp_1124;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1126 <= _tmp_1125;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1127 <= _tmp_1126;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1128 <= _tmp_1127;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1129 <= _tmp_1128;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1130 <= _tmp_1129;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1131 <= _tmp_1130;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1132 <= cparam_max_pool_47_stream_size;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1133 <= _tmp_1132;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1134 <= _tmp_1133;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1135 <= _tmp_1134;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1136 <= _tmp_1135;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1137 <= _tmp_1136;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1138 <= _tmp_1137;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1139 <= _tmp_1138;
      end 
      if(_tmp_1121) begin
        _stream_max_pool_47_sink_6_sink_mode <= 5'b1;
        _stream_max_pool_47_sink_6_sink_offset <= _tmp_1131;
        _stream_max_pool_47_sink_6_sink_size <= _tmp_1139;
        _stream_max_pool_47_sink_6_sink_stride <= 1;
      end 
      if(_tmp_1121) begin
        _stream_max_pool_47_sink_6_sink_sel <= 5;
      end 
      if(_stream_max_pool_47_sink_start && _stream_max_pool_47_sink_6_sink_mode & 5'b1 && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_sink_6_sink_offset_buf <= _stream_max_pool_47_sink_6_sink_offset;
        _stream_max_pool_47_sink_6_sink_size_buf <= _stream_max_pool_47_sink_6_sink_size;
        _stream_max_pool_47_sink_6_sink_stride_buf <= _stream_max_pool_47_sink_6_sink_stride;
      end 
      if((_stream_max_pool_47_sink_6_sink_fsm_4 == 1) && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_sink_6_sink_waddr <= _stream_max_pool_47_sink_6_sink_offset_buf - _stream_max_pool_47_sink_6_sink_stride_buf;
        _stream_max_pool_47_sink_6_sink_count <= _stream_max_pool_47_sink_6_sink_size_buf;
      end 
      if((_stream_max_pool_47_sink_6_sink_fsm_4 == 2) && _stream_max_pool_47_stream_oready) begin
        _stream_max_pool_47_sink_6_sink_waddr <= _stream_max_pool_47_sink_6_sink_waddr + _stream_max_pool_47_sink_6_sink_stride_buf;
        _stream_max_pool_47_sink_6_sink_wdata <= stream_max_pool_47_sink_6_data;
        _stream_max_pool_47_sink_6_sink_wenable <= 1;
        _stream_max_pool_47_sink_6_sink_count <= _stream_max_pool_47_sink_6_sink_count - 1;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1163 <= _stream_max_pool_47_source_start;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1164 <= _tmp_1163;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1165 <= _tmp_1164;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1168 <= _tmp_1167;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1169 <= _stream_max_pool_47_source_start;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1170 <= _tmp_1169;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1171 <= _tmp_1170;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1172 <= _tmp_1171;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1173 <= _tmp_1172;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1174 <= _tmp_1173;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1175 <= _tmp_1174;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1176 <= _tmp_1175;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1177 <= _stream_max_pool_47_source_stop;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1178 <= _tmp_1177;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1179 <= _tmp_1178;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1180 <= _tmp_1179;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1181 <= _tmp_1180;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1182 <= _tmp_1181;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1183 <= _tmp_1182;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1184 <= _tmp_1183;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1185 <= _stream_max_pool_47_source_busy;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1186 <= _tmp_1185;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1187 <= _tmp_1186;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1188 <= _tmp_1187;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1189 <= _tmp_1188;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1190 <= _tmp_1189;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1191 <= _tmp_1190;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1192 <= _tmp_1191;
      end 
      if(_stream_max_pool_47_stream_oready) begin
        _tmp_1193 <= _stream_max_pool_47_sink_busy;
      end 
      if(!_stream_max_pool_47_sink_busy && _tmp_1193) begin
        _stream_max_pool_47_busy_reg <= 0;
      end 
      if(_stream_max_pool_47_source_busy) begin
        _stream_max_pool_47_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_max_pool_47_fsm_1 = 1;
  localparam _stream_max_pool_47_fsm_2 = 2;
  localparam _stream_max_pool_47_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_47_fsm <= _stream_max_pool_47_fsm_init;
      _stream_max_pool_47_source_start <= 0;
      _stream_max_pool_47_source_busy <= 0;
      _stream_max_pool_47_stream_ivalid <= 0;
    end else begin
      if(_stream_max_pool_47_stream_oready && _tmp_1165) begin
        _stream_max_pool_47_stream_ivalid <= 1;
      end 
      if(_stream_max_pool_47_stream_oready && _tmp_1168) begin
        _stream_max_pool_47_stream_ivalid <= 0;
      end 
      case(_stream_max_pool_47_fsm)
        _stream_max_pool_47_fsm_init: begin
          if(_stream_max_pool_47_run_flag) begin
            _stream_max_pool_47_source_start <= 1;
          end 
          if(_stream_max_pool_47_run_flag) begin
            _stream_max_pool_47_fsm <= _stream_max_pool_47_fsm_1;
          end 
        end
        _stream_max_pool_47_fsm_1: begin
          if(_stream_max_pool_47_source_start && _stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_source_start <= 0;
            _stream_max_pool_47_source_busy <= 1;
          end 
          if(_stream_max_pool_47_source_start && _stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_fsm <= _stream_max_pool_47_fsm_2;
          end 
        end
        _stream_max_pool_47_fsm_2: begin
          if(_stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_fsm <= _stream_max_pool_47_fsm_3;
          end 
        end
        _stream_max_pool_47_fsm_3: begin
          if(_stream_max_pool_47_stream_oready && (_stream_max_pool_47_source_1_idle && _stream_max_pool_47_source_2_idle && _stream_max_pool_47_source_3_idle && _stream_max_pool_47_source_4_idle && (_stream_max_pool_47_fsm == 3))) begin
            _stream_max_pool_47_source_busy <= 0;
          end 
          if(_stream_max_pool_47_stream_oready && (_stream_max_pool_47_source_1_idle && _stream_max_pool_47_source_2_idle && _stream_max_pool_47_source_3_idle && _stream_max_pool_47_source_4_idle && (_stream_max_pool_47_fsm == 3)) && _stream_max_pool_47_run_flag) begin
            _stream_max_pool_47_source_start <= 1;
          end 
          if(_stream_max_pool_47_stream_oready && (_stream_max_pool_47_source_1_idle && _stream_max_pool_47_source_2_idle && _stream_max_pool_47_source_3_idle && _stream_max_pool_47_source_4_idle && (_stream_max_pool_47_fsm == 3))) begin
            _stream_max_pool_47_fsm <= _stream_max_pool_47_fsm_init;
          end 
          if(_stream_max_pool_47_stream_oready && (_stream_max_pool_47_source_1_idle && _stream_max_pool_47_source_2_idle && _stream_max_pool_47_source_3_idle && _stream_max_pool_47_source_4_idle && (_stream_max_pool_47_fsm == 3)) && _stream_max_pool_47_run_flag) begin
            _stream_max_pool_47_fsm <= _stream_max_pool_47_fsm_1;
          end 
        end
      endcase
    end
  end

  localparam main_fsm_1 = 1;
  localparam main_fsm_2 = 2;
  localparam main_fsm_3 = 3;
  localparam main_fsm_4 = 4;
  localparam main_fsm_5 = 5;
  localparam main_fsm_6 = 6;
  localparam main_fsm_7 = 7;
  localparam main_fsm_8 = 8;
  localparam main_fsm_9 = 9;
  localparam main_fsm_10 = 10;
  localparam main_fsm_11 = 11;
  localparam main_fsm_12 = 12;
  localparam main_fsm_13 = 13;
  localparam main_fsm_14 = 14;
  localparam main_fsm_15 = 15;
  localparam main_fsm_16 = 16;
  localparam main_fsm_17 = 17;
  localparam main_fsm_18 = 18;
  localparam main_fsm_19 = 19;
  localparam main_fsm_20 = 20;
  localparam main_fsm_21 = 21;
  localparam main_fsm_22 = 22;
  localparam main_fsm_23 = 23;
  localparam main_fsm_24 = 24;
  localparam main_fsm_25 = 25;
  localparam main_fsm_26 = 26;
  localparam main_fsm_27 = 27;
  localparam main_fsm_28 = 28;
  localparam main_fsm_29 = 29;
  localparam main_fsm_30 = 30;
  localparam main_fsm_31 = 31;
  localparam main_fsm_32 = 32;
  localparam main_fsm_33 = 33;
  localparam main_fsm_34 = 34;
  localparam main_fsm_35 = 35;
  localparam main_fsm_36 = 36;
  localparam main_fsm_37 = 37;
  localparam main_fsm_38 = 38;
  localparam main_fsm_39 = 39;
  localparam main_fsm_40 = 40;
  localparam main_fsm_41 = 41;
  localparam main_fsm_42 = 42;
  localparam main_fsm_43 = 43;
  localparam main_fsm_44 = 44;
  localparam main_fsm_45 = 45;
  localparam main_fsm_46 = 46;
  localparam main_fsm_47 = 47;
  localparam main_fsm_48 = 48;
  localparam main_fsm_49 = 49;
  localparam main_fsm_50 = 50;
  localparam main_fsm_51 = 51;
  localparam main_fsm_52 = 52;
  localparam main_fsm_53 = 53;
  localparam main_fsm_54 = 54;
  localparam main_fsm_55 = 55;
  localparam main_fsm_56 = 56;
  localparam main_fsm_57 = 57;
  localparam main_fsm_58 = 58;
  localparam main_fsm_59 = 59;
  localparam main_fsm_60 = 60;
  localparam main_fsm_61 = 61;
  localparam main_fsm_62 = 62;
  localparam main_fsm_63 = 63;
  localparam main_fsm_64 = 64;
  localparam main_fsm_65 = 65;
  localparam main_fsm_66 = 66;
  localparam main_fsm_67 = 67;
  localparam main_fsm_68 = 68;
  localparam main_fsm_69 = 69;
  localparam main_fsm_70 = 70;
  localparam main_fsm_71 = 71;
  localparam main_fsm_72 = 72;
  localparam main_fsm_73 = 73;
  localparam main_fsm_74 = 74;
  localparam main_fsm_75 = 75;
  localparam main_fsm_76 = 76;
  localparam main_fsm_77 = 77;
  localparam main_fsm_78 = 78;
  localparam main_fsm_79 = 79;
  localparam main_fsm_80 = 80;
  localparam main_fsm_81 = 81;
  localparam main_fsm_82 = 82;
  localparam main_fsm_83 = 83;
  localparam main_fsm_84 = 84;
  localparam main_fsm_85 = 85;
  localparam main_fsm_86 = 86;
  localparam main_fsm_87 = 87;
  localparam main_fsm_88 = 88;
  localparam main_fsm_89 = 89;
  localparam main_fsm_90 = 90;
  localparam main_fsm_91 = 91;
  localparam main_fsm_92 = 92;
  localparam main_fsm_93 = 93;
  localparam main_fsm_94 = 94;
  localparam main_fsm_95 = 95;
  localparam main_fsm_96 = 96;
  localparam main_fsm_97 = 97;
  localparam main_fsm_98 = 98;
  localparam main_fsm_99 = 99;
  localparam main_fsm_100 = 100;
  localparam main_fsm_101 = 101;
  localparam main_fsm_102 = 102;
  localparam main_fsm_103 = 103;
  localparam main_fsm_104 = 104;
  localparam main_fsm_105 = 105;
  localparam main_fsm_106 = 106;
  localparam main_fsm_107 = 107;
  localparam main_fsm_108 = 108;
  localparam main_fsm_109 = 109;
  localparam main_fsm_110 = 110;
  localparam main_fsm_111 = 111;
  localparam main_fsm_112 = 112;
  localparam main_fsm_113 = 113;
  localparam main_fsm_114 = 114;
  localparam main_fsm_115 = 115;
  localparam main_fsm_116 = 116;
  localparam main_fsm_117 = 117;
  localparam main_fsm_118 = 118;
  localparam main_fsm_119 = 119;
  localparam main_fsm_120 = 120;

  always @(posedge CLK) begin
    if(RST) begin
      main_fsm <= main_fsm_init;
      conv2d_25_objaddr <= 0;
      conv2d_25_arg_objaddr_0 <= 0;
      conv2d_25_arg_objaddr_1 <= 0;
      conv2d_25_arg_objaddr_2 <= 0;
      conv2d_25_arg_objaddr_3 <= 0;
      conv2d_25_control_param_index <= 0;
      max_pool_serial_27_objaddr <= 0;
      max_pool_serial_27_arg_objaddr_0 <= 0;
      max_pool_serial_27_control_param_index <= 0;
      max_pool_47_objaddr <= 0;
      max_pool_47_arg_objaddr_0 <= 0;
    end else begin
      case(main_fsm)
        main_fsm_init: begin
          if(_saxi_register_4 != 0) begin
            main_fsm <= main_fsm_1;
          end 
        end
        main_fsm_1: begin
          main_fsm <= main_fsm_2;
        end
        main_fsm_2: begin
          main_fsm <= main_fsm_3;
        end
        main_fsm_3: begin
          main_fsm <= main_fsm_4;
        end
        main_fsm_4: begin
          main_fsm <= main_fsm_5;
        end
        main_fsm_5: begin
          conv2d_25_objaddr <= _saxi_register_33;
          main_fsm <= main_fsm_6;
        end
        main_fsm_6: begin
          conv2d_25_arg_objaddr_0 <= _saxi_register_35;
          main_fsm <= main_fsm_7;
        end
        main_fsm_7: begin
          conv2d_25_arg_objaddr_1 <= _saxi_register_36;
          main_fsm <= main_fsm_8;
        end
        main_fsm_8: begin
          conv2d_25_arg_objaddr_2 <= _saxi_register_36 + 1728;
          main_fsm <= main_fsm_9;
        end
        main_fsm_9: begin
          conv2d_25_arg_objaddr_3 <= _saxi_register_36 + 1792;
          main_fsm <= main_fsm_10;
        end
        main_fsm_10: begin
          conv2d_25_control_param_index <= 0;
          main_fsm <= main_fsm_11;
        end
        main_fsm_11: begin
          main_fsm <= main_fsm_12;
        end
        main_fsm_12: begin
          main_fsm <= main_fsm_13;
        end
        main_fsm_13: begin
          if(control_conv2d_25 == 34) begin
            main_fsm <= main_fsm_14;
          end 
        end
        main_fsm_14: begin
          main_fsm <= main_fsm_15;
        end
        main_fsm_15: begin
          max_pool_serial_27_objaddr <= _saxi_register_33 + 11075584;
          main_fsm <= main_fsm_16;
        end
        main_fsm_16: begin
          max_pool_serial_27_arg_objaddr_0 <= _saxi_register_33;
          main_fsm <= main_fsm_17;
        end
        main_fsm_17: begin
          max_pool_serial_27_control_param_index <= 0;
          main_fsm <= main_fsm_18;
        end
        main_fsm_18: begin
          main_fsm <= main_fsm_19;
        end
        main_fsm_19: begin
          main_fsm <= main_fsm_20;
        end
        main_fsm_20: begin
          if(control_max_pool_serial_27 == 19) begin
            main_fsm <= main_fsm_21;
          end 
        end
        main_fsm_21: begin
          main_fsm <= main_fsm_22;
        end
        main_fsm_22: begin
          conv2d_25_objaddr <= _saxi_register_33 + 13844480;
          main_fsm <= main_fsm_23;
        end
        main_fsm_23: begin
          conv2d_25_arg_objaddr_0 <= _saxi_register_33 + 11075584;
          main_fsm <= main_fsm_24;
        end
        main_fsm_24: begin
          conv2d_25_arg_objaddr_1 <= _saxi_register_36 + 1856;
          main_fsm <= main_fsm_25;
        end
        main_fsm_25: begin
          conv2d_25_arg_objaddr_2 <= _saxi_register_36 + 20288;
          main_fsm <= main_fsm_26;
        end
        main_fsm_26: begin
          conv2d_25_arg_objaddr_3 <= _saxi_register_36 + 20416;
          main_fsm <= main_fsm_27;
        end
        main_fsm_27: begin
          conv2d_25_control_param_index <= 1;
          main_fsm <= main_fsm_28;
        end
        main_fsm_28: begin
          main_fsm <= main_fsm_29;
        end
        main_fsm_29: begin
          main_fsm <= main_fsm_30;
        end
        main_fsm_30: begin
          if(control_conv2d_25 == 34) begin
            main_fsm <= main_fsm_31;
          end 
        end
        main_fsm_31: begin
          main_fsm <= main_fsm_32;
        end
        main_fsm_32: begin
          max_pool_serial_27_objaddr <= _saxi_register_33 + 19382272;
          main_fsm <= main_fsm_33;
        end
        main_fsm_33: begin
          max_pool_serial_27_arg_objaddr_0 <= _saxi_register_33 + 13844480;
          main_fsm <= main_fsm_34;
        end
        main_fsm_34: begin
          max_pool_serial_27_control_param_index <= 1;
          main_fsm <= main_fsm_35;
        end
        main_fsm_35: begin
          main_fsm <= main_fsm_36;
        end
        main_fsm_36: begin
          main_fsm <= main_fsm_37;
        end
        main_fsm_37: begin
          if(control_max_pool_serial_27 == 19) begin
            main_fsm <= main_fsm_38;
          end 
        end
        main_fsm_38: begin
          main_fsm <= main_fsm_39;
        end
        main_fsm_39: begin
          conv2d_25_objaddr <= _saxi_register_33 + 20766720;
          main_fsm <= main_fsm_40;
        end
        main_fsm_40: begin
          conv2d_25_arg_objaddr_0 <= _saxi_register_33 + 19382272;
          main_fsm <= main_fsm_41;
        end
        main_fsm_41: begin
          conv2d_25_arg_objaddr_1 <= _saxi_register_36 + 20480;
          main_fsm <= main_fsm_42;
        end
        main_fsm_42: begin
          conv2d_25_arg_objaddr_2 <= _saxi_register_36 + 94208;
          main_fsm <= main_fsm_43;
        end
        main_fsm_43: begin
          conv2d_25_arg_objaddr_3 <= _saxi_register_36 + 94464;
          main_fsm <= main_fsm_44;
        end
        main_fsm_44: begin
          conv2d_25_control_param_index <= 2;
          main_fsm <= main_fsm_45;
        end
        main_fsm_45: begin
          main_fsm <= main_fsm_46;
        end
        main_fsm_46: begin
          main_fsm <= main_fsm_47;
        end
        main_fsm_47: begin
          if(control_conv2d_25 == 34) begin
            main_fsm <= main_fsm_48;
          end 
        end
        main_fsm_48: begin
          main_fsm <= main_fsm_49;
        end
        main_fsm_49: begin
          max_pool_serial_27_objaddr <= _saxi_register_33 + 23535616;
          main_fsm <= main_fsm_50;
        end
        main_fsm_50: begin
          max_pool_serial_27_arg_objaddr_0 <= _saxi_register_33 + 20766720;
          main_fsm <= main_fsm_51;
        end
        main_fsm_51: begin
          max_pool_serial_27_control_param_index <= 2;
          main_fsm <= main_fsm_52;
        end
        main_fsm_52: begin
          main_fsm <= main_fsm_53;
        end
        main_fsm_53: begin
          main_fsm <= main_fsm_54;
        end
        main_fsm_54: begin
          if(control_max_pool_serial_27 == 19) begin
            main_fsm <= main_fsm_55;
          end 
        end
        main_fsm_55: begin
          main_fsm <= main_fsm_56;
        end
        main_fsm_56: begin
          conv2d_25_objaddr <= _saxi_register_33 + 24227840;
          main_fsm <= main_fsm_57;
        end
        main_fsm_57: begin
          conv2d_25_arg_objaddr_0 <= _saxi_register_33 + 23535616;
          main_fsm <= main_fsm_58;
        end
        main_fsm_58: begin
          conv2d_25_arg_objaddr_1 <= _saxi_register_36 + 94528;
          main_fsm <= main_fsm_59;
        end
        main_fsm_59: begin
          conv2d_25_arg_objaddr_2 <= _saxi_register_36 + 389440;
          main_fsm <= main_fsm_60;
        end
        main_fsm_60: begin
          conv2d_25_arg_objaddr_3 <= _saxi_register_36 + 389952;
          main_fsm <= main_fsm_61;
        end
        main_fsm_61: begin
          conv2d_25_control_param_index <= 3;
          main_fsm <= main_fsm_62;
        end
        main_fsm_62: begin
          main_fsm <= main_fsm_63;
        end
        main_fsm_63: begin
          main_fsm <= main_fsm_64;
        end
        main_fsm_64: begin
          if(control_conv2d_25 == 34) begin
            main_fsm <= main_fsm_65;
          end 
        end
        main_fsm_65: begin
          main_fsm <= main_fsm_66;
        end
        main_fsm_66: begin
          max_pool_serial_27_objaddr <= _saxi_register_33 + 25612288;
          main_fsm <= main_fsm_67;
        end
        main_fsm_67: begin
          max_pool_serial_27_arg_objaddr_0 <= _saxi_register_33 + 24227840;
          main_fsm <= main_fsm_68;
        end
        main_fsm_68: begin
          max_pool_serial_27_control_param_index <= 3;
          main_fsm <= main_fsm_69;
        end
        main_fsm_69: begin
          main_fsm <= main_fsm_70;
        end
        main_fsm_70: begin
          main_fsm <= main_fsm_71;
        end
        main_fsm_71: begin
          if(control_max_pool_serial_27 == 19) begin
            main_fsm <= main_fsm_72;
          end 
        end
        main_fsm_72: begin
          main_fsm <= main_fsm_73;
        end
        main_fsm_73: begin
          conv2d_25_objaddr <= _saxi_register_33 + 25958400;
          main_fsm <= main_fsm_74;
        end
        main_fsm_74: begin
          conv2d_25_arg_objaddr_0 <= _saxi_register_33 + 25612288;
          main_fsm <= main_fsm_75;
        end
        main_fsm_75: begin
          conv2d_25_arg_objaddr_1 <= _saxi_register_36 + 390016;
          main_fsm <= main_fsm_76;
        end
        main_fsm_76: begin
          conv2d_25_arg_objaddr_2 <= _saxi_register_36 + 1569664;
          main_fsm <= main_fsm_77;
        end
        main_fsm_77: begin
          conv2d_25_arg_objaddr_3 <= _saxi_register_36 + 1570688;
          main_fsm <= main_fsm_78;
        end
        main_fsm_78: begin
          conv2d_25_control_param_index <= 4;
          main_fsm <= main_fsm_79;
        end
        main_fsm_79: begin
          main_fsm <= main_fsm_80;
        end
        main_fsm_80: begin
          main_fsm <= main_fsm_81;
        end
        main_fsm_81: begin
          if(control_conv2d_25 == 34) begin
            main_fsm <= main_fsm_82;
          end 
        end
        main_fsm_82: begin
          main_fsm <= main_fsm_83;
        end
        main_fsm_83: begin
          max_pool_serial_27_objaddr <= _saxi_register_33 + 26650624;
          main_fsm <= main_fsm_84;
        end
        main_fsm_84: begin
          max_pool_serial_27_arg_objaddr_0 <= _saxi_register_33 + 25958400;
          main_fsm <= main_fsm_85;
        end
        main_fsm_85: begin
          max_pool_serial_27_control_param_index <= 4;
          main_fsm <= main_fsm_86;
        end
        main_fsm_86: begin
          main_fsm <= main_fsm_87;
        end
        main_fsm_87: begin
          main_fsm <= main_fsm_88;
        end
        main_fsm_88: begin
          if(control_max_pool_serial_27 == 19) begin
            main_fsm <= main_fsm_89;
          end 
        end
        main_fsm_89: begin
          main_fsm <= main_fsm_90;
        end
        main_fsm_90: begin
          conv2d_25_objaddr <= _saxi_register_33 + 26823680;
          main_fsm <= main_fsm_91;
        end
        main_fsm_91: begin
          conv2d_25_arg_objaddr_0 <= _saxi_register_33 + 26650624;
          main_fsm <= main_fsm_92;
        end
        main_fsm_92: begin
          conv2d_25_arg_objaddr_1 <= _saxi_register_36 + 1570752;
          main_fsm <= main_fsm_93;
        end
        main_fsm_93: begin
          conv2d_25_arg_objaddr_2 <= _saxi_register_36 + 6289344;
          main_fsm <= main_fsm_94;
        end
        main_fsm_94: begin
          conv2d_25_arg_objaddr_3 <= _saxi_register_36 + 6291392;
          main_fsm <= main_fsm_95;
        end
        main_fsm_95: begin
          conv2d_25_control_param_index <= 5;
          main_fsm <= main_fsm_96;
        end
        main_fsm_96: begin
          main_fsm <= main_fsm_97;
        end
        main_fsm_97: begin
          main_fsm <= main_fsm_98;
        end
        main_fsm_98: begin
          if(control_conv2d_25 == 34) begin
            main_fsm <= main_fsm_99;
          end 
        end
        main_fsm_99: begin
          main_fsm <= main_fsm_100;
        end
        main_fsm_100: begin
          max_pool_47_objaddr <= _saxi_register_33 + 27169792;
          main_fsm <= main_fsm_101;
        end
        main_fsm_101: begin
          max_pool_47_arg_objaddr_0 <= _saxi_register_33 + 26823680;
          main_fsm <= main_fsm_102;
        end
        main_fsm_102: begin
          main_fsm <= main_fsm_103;
        end
        main_fsm_103: begin
          main_fsm <= main_fsm_104;
        end
        main_fsm_104: begin
          if(control_max_pool_47 == 19) begin
            main_fsm <= main_fsm_105;
          end 
        end
        main_fsm_105: begin
          main_fsm <= main_fsm_106;
        end
        main_fsm_106: begin
          conv2d_25_objaddr <= _saxi_register_34;
          main_fsm <= main_fsm_107;
        end
        main_fsm_107: begin
          conv2d_25_arg_objaddr_0 <= _saxi_register_33 + 27169792;
          main_fsm <= main_fsm_108;
        end
        main_fsm_108: begin
          conv2d_25_arg_objaddr_1 <= _saxi_register_36 + 6291456;
          main_fsm <= main_fsm_109;
        end
        main_fsm_109: begin
          conv2d_25_arg_objaddr_2 <= _saxi_register_36 + 25165824;
          main_fsm <= main_fsm_110;
        end
        main_fsm_110: begin
          conv2d_25_arg_objaddr_3 <= _saxi_register_36 + 25169920;
          main_fsm <= main_fsm_111;
        end
        main_fsm_111: begin
          conv2d_25_control_param_index <= 6;
          main_fsm <= main_fsm_112;
        end
        main_fsm_112: begin
          main_fsm <= main_fsm_113;
        end
        main_fsm_113: begin
          main_fsm <= main_fsm_114;
        end
        main_fsm_114: begin
          if(control_conv2d_25 == 34) begin
            main_fsm <= main_fsm_115;
          end 
        end
        main_fsm_115: begin
          main_fsm <= main_fsm_116;
        end
        main_fsm_116: begin
          main_fsm <= main_fsm_117;
        end
        main_fsm_117: begin
          main_fsm <= main_fsm_118;
        end
        main_fsm_118: begin
          main_fsm <= main_fsm_119;
        end
        main_fsm_119: begin
          main_fsm <= main_fsm_120;
        end
        main_fsm_120: begin
          main_fsm <= main_fsm_init;
        end
      endcase
    end
  end

  localparam control_conv2d_25_1 = 1;
  localparam control_conv2d_25_2 = 2;
  localparam control_conv2d_25_3 = 3;
  localparam control_conv2d_25_4 = 4;
  localparam control_conv2d_25_5 = 5;
  localparam control_conv2d_25_6 = 6;
  localparam control_conv2d_25_7 = 7;
  localparam control_conv2d_25_8 = 8;
  localparam control_conv2d_25_9 = 9;
  localparam control_conv2d_25_10 = 10;
  localparam control_conv2d_25_11 = 11;
  localparam control_conv2d_25_12 = 12;
  localparam control_conv2d_25_13 = 13;
  localparam control_conv2d_25_14 = 14;
  localparam control_conv2d_25_15 = 15;
  localparam control_conv2d_25_16 = 16;
  localparam control_conv2d_25_17 = 17;
  localparam control_conv2d_25_18 = 18;
  localparam control_conv2d_25_19 = 19;
  localparam control_conv2d_25_20 = 20;
  localparam control_conv2d_25_21 = 21;
  localparam control_conv2d_25_22 = 22;
  localparam control_conv2d_25_23 = 23;
  localparam control_conv2d_25_24 = 24;
  localparam control_conv2d_25_25 = 25;
  localparam control_conv2d_25_26 = 26;
  localparam control_conv2d_25_27 = 27;
  localparam control_conv2d_25_28 = 28;
  localparam control_conv2d_25_29 = 29;
  localparam control_conv2d_25_30 = 30;
  localparam control_conv2d_25_31 = 31;
  localparam control_conv2d_25_32 = 32;
  localparam control_conv2d_25_33 = 33;
  localparam control_conv2d_25_34 = 34;

  always @(posedge CLK) begin
    if(RST) begin
      control_conv2d_25 <= control_conv2d_25_init;
      _control_conv2d_25_called <= 0;
      conv2d_25_filter_base_offset <= 0;
      conv2d_25_filter_page_comp_offset <= 0;
      conv2d_25_filter_page_dma_offset <= 0;
      conv2d_25_act_base_offset_row <= 0;
      conv2d_25_act_base_offset_bat <= 0;
      conv2d_25_dma_flag_0 <= 0;
      conv2d_25_dma_flag_1 <= 0;
      conv2d_25_dma_flag_2 <= 0;
      conv2d_25_act_page_comp_offset_0 <= 0;
      conv2d_25_act_page_comp_offset_1 <= 0;
      conv2d_25_act_page_comp_offset_2 <= 0;
      conv2d_25_act_page_dma_offset_0 <= 0;
      conv2d_25_act_page_dma_offset_1 <= 0;
      conv2d_25_act_page_dma_offset_2 <= 0;
      conv2d_25_out_base_offset_val <= 0;
      conv2d_25_out_base_offset_col <= 0;
      conv2d_25_out_base_offset_row <= 0;
      conv2d_25_out_base_offset_bat <= 0;
      conv2d_25_out_base_offset_och <= 0;
      conv2d_25_out_page <= 0;
      conv2d_25_out_page_comp_offset <= 0;
      conv2d_25_out_page_dma_offset <= 0;
      conv2d_25_out_laddr_offset <= 0;
      conv2d_25_sync_out_count <= 0;
      conv2d_25_write_count <= 0;
      conv2d_25_next_out_write_size <= 0;
      conv2d_25_row_count <= 0;
      conv2d_25_bat_count <= 0;
      conv2d_25_och_count <= 0;
      conv2d_25_row_select <= 0;
      conv2d_25_prev_row_count <= 0;
      conv2d_25_prev_bat_count <= 0;
      conv2d_25_prev_och_count <= 0;
      conv2d_25_prev_row_select <= 0;
      conv2d_25_out_col_count <= 0;
      conv2d_25_out_row_count <= 0;
      conv2d_25_out_ram_select <= 0;
      conv2d_25_skip_read_filter <= 0;
      conv2d_25_skip_read_act <= 0;
      conv2d_25_skip_comp <= 0;
      conv2d_25_skip_write_out <= 1;
    end else begin
      case(control_conv2d_25)
        control_conv2d_25_init: begin
          if(main_fsm == 11) begin
            _control_conv2d_25_called <= 1;
          end 
          if(main_fsm == 28) begin
            _control_conv2d_25_called <= 1;
          end 
          if(main_fsm == 45) begin
            _control_conv2d_25_called <= 1;
          end 
          if(main_fsm == 62) begin
            _control_conv2d_25_called <= 1;
          end 
          if(main_fsm == 79) begin
            _control_conv2d_25_called <= 1;
          end 
          if(main_fsm == 96) begin
            _control_conv2d_25_called <= 1;
          end 
          if(main_fsm == 112) begin
            _control_conv2d_25_called <= 1;
          end 
          if(main_fsm == 11) begin
            control_conv2d_25 <= control_conv2d_25_1;
          end 
          if(main_fsm == 28) begin
            control_conv2d_25 <= control_conv2d_25_1;
          end 
          if(main_fsm == 45) begin
            control_conv2d_25 <= control_conv2d_25_1;
          end 
          if(main_fsm == 62) begin
            control_conv2d_25 <= control_conv2d_25_1;
          end 
          if(main_fsm == 79) begin
            control_conv2d_25 <= control_conv2d_25_1;
          end 
          if(main_fsm == 96) begin
            control_conv2d_25 <= control_conv2d_25_1;
          end 
          if(main_fsm == 112) begin
            control_conv2d_25 <= control_conv2d_25_1;
          end 
        end
        control_conv2d_25_1: begin
          control_conv2d_25 <= control_conv2d_25_2;
        end
        control_conv2d_25_2: begin
          conv2d_25_filter_base_offset <= 0;
          conv2d_25_filter_page_comp_offset <= 0;
          conv2d_25_filter_page_dma_offset <= 0;
          conv2d_25_act_base_offset_row <= 0;
          conv2d_25_act_base_offset_bat <= 0;
          conv2d_25_dma_flag_0 <= 1;
          conv2d_25_dma_flag_1 <= 1;
          conv2d_25_dma_flag_2 <= 1;
          conv2d_25_act_page_comp_offset_0 <= 0;
          conv2d_25_act_page_comp_offset_1 <= 0;
          conv2d_25_act_page_comp_offset_2 <= 0;
          conv2d_25_act_page_dma_offset_0 <= 0;
          conv2d_25_act_page_dma_offset_1 <= 0;
          conv2d_25_act_page_dma_offset_2 <= 0;
          conv2d_25_out_base_offset_val <= 0;
          conv2d_25_out_base_offset_col <= 0;
          conv2d_25_out_base_offset_row <= 0;
          conv2d_25_out_base_offset_bat <= 0;
          conv2d_25_out_base_offset_och <= 0;
          conv2d_25_out_page <= 0;
          conv2d_25_out_page_comp_offset <= 0;
          conv2d_25_out_page_dma_offset <= 0;
          conv2d_25_out_laddr_offset <= 0;
          conv2d_25_sync_out_count <= 0;
          conv2d_25_write_count <= 0;
          conv2d_25_next_out_write_size <= (cparam_conv2d_25_max_och_count == 0)? cparam_conv2d_25_out_write_size_res : cparam_conv2d_25_out_write_size;
          conv2d_25_row_count <= 0;
          conv2d_25_bat_count <= 0;
          conv2d_25_och_count <= 0;
          conv2d_25_row_select <= 0;
          conv2d_25_prev_row_count <= 0;
          conv2d_25_prev_bat_count <= 0;
          conv2d_25_prev_och_count <= 0;
          conv2d_25_prev_row_select <= 0;
          conv2d_25_out_col_count <= 0;
          conv2d_25_out_row_count <= 0;
          conv2d_25_out_ram_select <= 0;
          conv2d_25_skip_read_filter <= 0;
          conv2d_25_skip_read_act <= 0;
          conv2d_25_skip_comp <= 0;
          conv2d_25_skip_write_out <= 1;
          if(_maxi_read_req_idle) begin
            control_conv2d_25 <= control_conv2d_25_3;
          end 
        end
        control_conv2d_25_3: begin
          if(_maxi_read_idle) begin
            control_conv2d_25 <= control_conv2d_25_4;
          end 
        end
        control_conv2d_25_4: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_25 <= control_conv2d_25_5;
          end 
        end
        control_conv2d_25_5: begin
          if(_maxi_read_idle) begin
            control_conv2d_25 <= control_conv2d_25_6;
          end 
        end
        control_conv2d_25_6: begin
          if(cparam_conv2d_25_data_stationary == 0) begin
            control_conv2d_25 <= control_conv2d_25_7;
          end 
          if(cparam_conv2d_25_data_stationary == 1) begin
            control_conv2d_25 <= control_conv2d_25_12;
          end 
        end
        control_conv2d_25_7: begin
          control_conv2d_25 <= control_conv2d_25_8;
          if(conv2d_25_skip_read_filter) begin
            control_conv2d_25 <= control_conv2d_25_11;
          end 
        end
        control_conv2d_25_8: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_25 <= control_conv2d_25_9;
          end 
        end
        control_conv2d_25_9: begin
          if(_maxi_read_idle) begin
            control_conv2d_25 <= control_conv2d_25_10;
          end 
        end
        control_conv2d_25_10: begin
          control_conv2d_25 <= control_conv2d_25_11;
        end
        control_conv2d_25_11: begin
          if(cparam_conv2d_25_data_stationary == 0) begin
            control_conv2d_25 <= control_conv2d_25_12;
          end 
          if(cparam_conv2d_25_data_stationary == 1) begin
            control_conv2d_25 <= control_conv2d_25_24;
          end 
        end
        control_conv2d_25_12: begin
          control_conv2d_25 <= control_conv2d_25_13;
          if(conv2d_25_skip_read_act) begin
            control_conv2d_25 <= control_conv2d_25_23;
          end 
        end
        control_conv2d_25_13: begin
          control_conv2d_25 <= control_conv2d_25_14;
          if(conv2d_25_mux_dma_pad_mask_0 || !conv2d_25_mux_dma_flag_0) begin
            control_conv2d_25 <= control_conv2d_25_16;
          end 
        end
        control_conv2d_25_14: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_25 <= control_conv2d_25_15;
          end 
        end
        control_conv2d_25_15: begin
          if(_maxi_read_idle) begin
            control_conv2d_25 <= control_conv2d_25_16;
          end 
        end
        control_conv2d_25_16: begin
          control_conv2d_25 <= control_conv2d_25_17;
          if(conv2d_25_mux_dma_pad_mask_1 || !conv2d_25_mux_dma_flag_1) begin
            control_conv2d_25 <= control_conv2d_25_19;
          end 
        end
        control_conv2d_25_17: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_25 <= control_conv2d_25_18;
          end 
        end
        control_conv2d_25_18: begin
          if(_maxi_read_idle) begin
            control_conv2d_25 <= control_conv2d_25_19;
          end 
        end
        control_conv2d_25_19: begin
          control_conv2d_25 <= control_conv2d_25_20;
          if(conv2d_25_mux_dma_pad_mask_2 || !conv2d_25_mux_dma_flag_2) begin
            control_conv2d_25 <= control_conv2d_25_22;
          end 
        end
        control_conv2d_25_20: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_25 <= control_conv2d_25_21;
          end 
        end
        control_conv2d_25_21: begin
          if(_maxi_read_idle) begin
            control_conv2d_25 <= control_conv2d_25_22;
          end 
        end
        control_conv2d_25_22: begin
          control_conv2d_25 <= control_conv2d_25_23;
        end
        control_conv2d_25_23: begin
          if(cparam_conv2d_25_data_stationary == 0) begin
            control_conv2d_25 <= control_conv2d_25_24;
          end 
          if(cparam_conv2d_25_data_stationary == 1) begin
            control_conv2d_25 <= control_conv2d_25_7;
          end 
        end
        control_conv2d_25_24: begin
          if(_maxi_write_idle) begin
            control_conv2d_25 <= control_conv2d_25_25;
          end 
        end
        control_conv2d_25_25: begin
          if(conv2d_25_comp_fsm == 0) begin
            control_conv2d_25 <= control_conv2d_25_26;
          end 
        end
        control_conv2d_25_26: begin
          control_conv2d_25 <= control_conv2d_25_27;
          if(conv2d_25_skip_write_out) begin
            control_conv2d_25 <= control_conv2d_25_32;
          end 
          if((cparam_conv2d_25_data_stationary == 1) && (conv2d_25_prev_och_count < cparam_conv2d_25_max_och_count)) begin
            control_conv2d_25 <= control_conv2d_25_32;
          end 
        end
        control_conv2d_25_27: begin
          if(conv2d_25_sync_comp_count >= conv2d_25_sync_out_count + cparam_conv2d_25_inc_sync_out) begin
            control_conv2d_25 <= control_conv2d_25_28;
          end 
        end
        control_conv2d_25_28: begin
          if(!conv2d_25_dma_out_mask_0) begin
            control_conv2d_25 <= control_conv2d_25_29;
          end 
          if(conv2d_25_dma_out_mask_0) begin
            control_conv2d_25 <= control_conv2d_25_30;
          end 
        end
        control_conv2d_25_29: begin
          if(_maxi_write_req_idle) begin
            control_conv2d_25 <= control_conv2d_25_30;
          end 
        end
        control_conv2d_25_30: begin
          control_conv2d_25 <= control_conv2d_25_31;
        end
        control_conv2d_25_31: begin
          conv2d_25_write_count <= conv2d_25_write_count + 1;
          if(conv2d_25_out_ram_select == 0) begin
            conv2d_25_out_laddr_offset <= conv2d_25_out_laddr_offset + conv2d_25_next_out_write_size;
          end 
          if((cparam_conv2d_25_data_stationary == 0) && !cparam_conv2d_25_keep_filter) begin
            conv2d_25_out_base_offset_col <= conv2d_25_out_base_offset_col + cparam_conv2d_25_out_col_step;
            conv2d_25_out_col_count <= conv2d_25_out_col_count + 1;
          end 
          conv2d_25_out_ram_select <= conv2d_25_out_ram_select + 1;
          if(conv2d_25_out_ram_select == 0) begin
            conv2d_25_out_ram_select <= 0;
          end 
          conv2d_25_sync_out_count <= conv2d_25_sync_out_count + cparam_conv2d_25_inc_sync_out;
          if((cparam_conv2d_25_data_stationary == 0) && !cparam_conv2d_25_keep_filter && (conv2d_25_write_count >= cparam_conv2d_25_out_num_col - 1) || (cparam_conv2d_25_data_stationary == 0) && cparam_conv2d_25_keep_filter || (cparam_conv2d_25_data_stationary == 1)) begin
            conv2d_25_sync_out_count <= conv2d_25_sync_out_count + (cparam_conv2d_25_inc_sync_out + cparam_conv2d_25_inc_sync_out_res);
          end 
          if((cparam_conv2d_25_data_stationary == 0) && !cparam_conv2d_25_keep_filter) begin
            control_conv2d_25 <= control_conv2d_25_26;
          end 
          if((cparam_conv2d_25_data_stationary == 0) && !cparam_conv2d_25_keep_filter && (conv2d_25_write_count >= cparam_conv2d_25_out_num_col - 1) || (cparam_conv2d_25_data_stationary == 0) && cparam_conv2d_25_keep_filter || (cparam_conv2d_25_data_stationary == 1)) begin
            control_conv2d_25 <= control_conv2d_25_32;
          end 
        end
        control_conv2d_25_32: begin
          if(conv2d_25_update_filter) begin
            conv2d_25_filter_base_offset <= conv2d_25_filter_base_offset + cparam_conv2d_25_filter_base_step;
          end 
          if((cparam_conv2d_25_data_stationary == 1) && (conv2d_25_och_count >= cparam_conv2d_25_max_och_count)) begin
            conv2d_25_filter_base_offset <= 0;
          end 
          if(conv2d_25_update_filter) begin
            conv2d_25_och_count <= conv2d_25_och_count + cparam_conv2d_25_och_count_step;
          end 
          if((cparam_conv2d_25_data_stationary == 1) && (conv2d_25_och_count >= cparam_conv2d_25_max_och_count)) begin
            conv2d_25_och_count <= 0;
          end 
          if(conv2d_25_update_filter) begin
            conv2d_25_filter_page_comp_offset <= conv2d_25_filter_page_comp_offset + cparam_conv2d_25_filter_read_step;
            conv2d_25_filter_page_dma_offset <= conv2d_25_filter_page_dma_offset + cparam_conv2d_25_filter_read_step;
          end 
          if(conv2d_25_update_filter && (conv2d_25_filter_page_comp_offset + cparam_conv2d_25_filter_read_step + cparam_conv2d_25_filter_read_step > 1024)) begin
            conv2d_25_filter_page_comp_offset <= 0;
            conv2d_25_filter_page_dma_offset <= 0;
          end 
          if(conv2d_25_update_act) begin
            conv2d_25_act_base_offset_row <= conv2d_25_act_base_offset_row + cparam_conv2d_25_act_row_step;
          end 
          if(conv2d_25_update_act && (conv2d_25_row_count >= cparam_conv2d_25_max_row_count)) begin
            conv2d_25_act_base_offset_row <= 0;
            conv2d_25_act_base_offset_bat <= conv2d_25_act_base_offset_bat + cparam_conv2d_25_act_bat_step;
          end 
          if(conv2d_25_update_act && (conv2d_25_row_count >= cparam_conv2d_25_max_row_count) && (conv2d_25_bat_count >= cparam_conv2d_25_max_bat_count)) begin
            conv2d_25_act_base_offset_bat <= 0;
          end 
          if(!conv2d_25_update_act) begin
            conv2d_25_dma_flag_0 <= 0;
          end 
          if(conv2d_25_update_act) begin
            conv2d_25_dma_flag_0 <= cparam_conv2d_25_dma_flag_conds_0;
          end 
          if(conv2d_25_update_act && (conv2d_25_row_count >= cparam_conv2d_25_max_row_count)) begin
            conv2d_25_dma_flag_0 <= 1;
          end 
          if(!conv2d_25_update_act) begin
            conv2d_25_dma_flag_1 <= 0;
          end 
          if(conv2d_25_update_act) begin
            conv2d_25_dma_flag_1 <= cparam_conv2d_25_dma_flag_conds_1;
          end 
          if(conv2d_25_update_act && (conv2d_25_row_count >= cparam_conv2d_25_max_row_count)) begin
            conv2d_25_dma_flag_1 <= 1;
          end 
          if(!conv2d_25_update_act) begin
            conv2d_25_dma_flag_2 <= 0;
          end 
          if(conv2d_25_update_act) begin
            conv2d_25_dma_flag_2 <= cparam_conv2d_25_dma_flag_conds_2;
          end 
          if(conv2d_25_update_act && (conv2d_25_row_count >= cparam_conv2d_25_max_row_count)) begin
            conv2d_25_dma_flag_2 <= 1;
          end 
          if(conv2d_25_update_act) begin
            conv2d_25_row_count <= conv2d_25_row_count + cparam_conv2d_25_stride_row_par_row;
          end 
          if(conv2d_25_update_act && (conv2d_25_row_count >= cparam_conv2d_25_max_row_count)) begin
            conv2d_25_row_count <= 0;
            conv2d_25_bat_count <= conv2d_25_bat_count + 1;
          end 
          if(conv2d_25_update_act && (conv2d_25_row_count >= cparam_conv2d_25_max_row_count) && (conv2d_25_bat_count >= cparam_conv2d_25_max_bat_count)) begin
            conv2d_25_bat_count <= 0;
          end 
          if(conv2d_25_update_act && (cparam_conv2d_25_stride_row_par_row < 3)) begin
            conv2d_25_row_select <= conv2d_25_row_select + cparam_conv2d_25_stride_row_par_row;
            conv2d_25_prev_row_select <= conv2d_25_row_select;
          end 
          if(conv2d_25_update_act && (cparam_conv2d_25_stride_row_par_row < 3) && (conv2d_25_row_select + cparam_conv2d_25_stride_row_par_row >= 3)) begin
            conv2d_25_row_select <= conv2d_25_row_select - (3 - cparam_conv2d_25_stride_row_par_row);
            conv2d_25_prev_row_select <= conv2d_25_row_select;
          end 
          if(conv2d_25_update_act && !(cparam_conv2d_25_stride_row_par_row < 3)) begin
            conv2d_25_row_select <= 0;
            conv2d_25_prev_row_select <= 0;
          end 
          if(conv2d_25_update_act && (conv2d_25_row_count >= cparam_conv2d_25_max_row_count)) begin
            conv2d_25_row_select <= 0;
            conv2d_25_prev_row_select <= 0;
          end 
          if(conv2d_25_update_act && conv2d_25_mux_next_dma_flag_0) begin
            conv2d_25_act_page_comp_offset_0 <= conv2d_25_act_page_comp_offset_0 + cparam_conv2d_25_act_read_step;
            conv2d_25_act_page_dma_offset_0 <= conv2d_25_act_page_dma_offset_0 + cparam_conv2d_25_act_read_step;
          end 
          if(conv2d_25_update_act && conv2d_25_mux_next_dma_flag_0 && (conv2d_25_act_page_comp_offset_0 + cparam_conv2d_25_act_read_step + cparam_conv2d_25_act_read_step > 4096)) begin
            conv2d_25_act_page_comp_offset_0 <= 0;
            conv2d_25_act_page_dma_offset_0 <= 0;
          end 
          if((cparam_conv2d_25_data_stationary == 0) && (conv2d_25_row_count >= cparam_conv2d_25_max_row_count) && (conv2d_25_bat_count >= cparam_conv2d_25_max_bat_count) && cparam_conv2d_25_keep_input) begin
            conv2d_25_act_page_comp_offset_0 <= 0;
            conv2d_25_act_page_dma_offset_0 <= 0;
          end 
          if(conv2d_25_update_act && conv2d_25_mux_next_dma_flag_1) begin
            conv2d_25_act_page_comp_offset_1 <= conv2d_25_act_page_comp_offset_1 + cparam_conv2d_25_act_read_step;
            conv2d_25_act_page_dma_offset_1 <= conv2d_25_act_page_dma_offset_1 + cparam_conv2d_25_act_read_step;
          end 
          if(conv2d_25_update_act && conv2d_25_mux_next_dma_flag_1 && (conv2d_25_act_page_comp_offset_1 + cparam_conv2d_25_act_read_step + cparam_conv2d_25_act_read_step > 4096)) begin
            conv2d_25_act_page_comp_offset_1 <= 0;
            conv2d_25_act_page_dma_offset_1 <= 0;
          end 
          if((cparam_conv2d_25_data_stationary == 0) && (conv2d_25_row_count >= cparam_conv2d_25_max_row_count) && (conv2d_25_bat_count >= cparam_conv2d_25_max_bat_count) && cparam_conv2d_25_keep_input) begin
            conv2d_25_act_page_comp_offset_1 <= 0;
            conv2d_25_act_page_dma_offset_1 <= 0;
          end 
          if(conv2d_25_update_act && conv2d_25_mux_next_dma_flag_2) begin
            conv2d_25_act_page_comp_offset_2 <= conv2d_25_act_page_comp_offset_2 + cparam_conv2d_25_act_read_step;
            conv2d_25_act_page_dma_offset_2 <= conv2d_25_act_page_dma_offset_2 + cparam_conv2d_25_act_read_step;
          end 
          if(conv2d_25_update_act && conv2d_25_mux_next_dma_flag_2 && (conv2d_25_act_page_comp_offset_2 + cparam_conv2d_25_act_read_step + cparam_conv2d_25_act_read_step > 4096)) begin
            conv2d_25_act_page_comp_offset_2 <= 0;
            conv2d_25_act_page_dma_offset_2 <= 0;
          end 
          if((cparam_conv2d_25_data_stationary == 0) && (conv2d_25_row_count >= cparam_conv2d_25_max_row_count) && (conv2d_25_bat_count >= cparam_conv2d_25_max_bat_count) && cparam_conv2d_25_keep_input) begin
            conv2d_25_act_page_comp_offset_2 <= 0;
            conv2d_25_act_page_dma_offset_2 <= 0;
          end 
          conv2d_25_next_out_write_size <= (conv2d_25_och_count >= cparam_conv2d_25_max_och_count)? cparam_conv2d_25_out_write_size_res : cparam_conv2d_25_out_write_size;
          if(!conv2d_25_skip_write_out) begin
            conv2d_25_write_count <= 0;
            conv2d_25_out_laddr_offset <= 0;
            conv2d_25_out_ram_select <= 0;
          end 
          if((cparam_conv2d_25_data_stationary == 0) && !conv2d_25_skip_write_out) begin
            conv2d_25_out_base_offset_col <= 0;
            conv2d_25_out_base_offset_row <= conv2d_25_out_base_offset_row + cparam_conv2d_25_out_row_step;
            conv2d_25_out_col_count <= 0;
            conv2d_25_out_row_count <= conv2d_25_out_row_count + 1;
          end 
          if((cparam_conv2d_25_data_stationary == 0) && !conv2d_25_skip_write_out && (conv2d_25_prev_row_count >= cparam_conv2d_25_max_row_count)) begin
            conv2d_25_out_base_offset_row <= 0;
            conv2d_25_out_base_offset_bat <= conv2d_25_out_base_offset_bat + cparam_conv2d_25_out_bat_step;
            conv2d_25_out_row_count <= 0;
          end 
          if((cparam_conv2d_25_data_stationary == 0) && !conv2d_25_skip_write_out && (conv2d_25_prev_row_count >= cparam_conv2d_25_max_row_count) && (conv2d_25_prev_bat_count >= cparam_conv2d_25_max_bat_count)) begin
            conv2d_25_out_base_offset_bat <= 0;
            conv2d_25_out_base_offset_och <= conv2d_25_out_base_offset_och + cparam_conv2d_25_out_och_step;
          end 
          if((cparam_conv2d_25_data_stationary == 1) && (conv2d_25_prev_och_count >= cparam_conv2d_25_max_och_count) && !conv2d_25_skip_write_out) begin
            conv2d_25_out_base_offset_row <= conv2d_25_out_base_offset_row + cparam_conv2d_25_out_row_step;
          end 
          if((cparam_conv2d_25_data_stationary == 0) && !conv2d_25_out_page) begin
            conv2d_25_out_page_comp_offset <= 512;
            conv2d_25_out_page_dma_offset <= 0;
            conv2d_25_out_page <= 1;
          end 
          if((cparam_conv2d_25_data_stationary == 0) && conv2d_25_out_page) begin
            conv2d_25_out_page_comp_offset <= 0;
            conv2d_25_out_page_dma_offset <= 512;
            conv2d_25_out_page <= 0;
          end 
          if((cparam_conv2d_25_data_stationary == 1) && (conv2d_25_och_count >= cparam_conv2d_25_max_och_count) && !conv2d_25_out_page) begin
            conv2d_25_out_page_comp_offset <= 512;
            conv2d_25_out_page_dma_offset <= 0;
            conv2d_25_out_page <= 1;
          end 
          if((cparam_conv2d_25_data_stationary == 1) && (conv2d_25_och_count >= cparam_conv2d_25_max_och_count) && conv2d_25_out_page) begin
            conv2d_25_out_page_comp_offset <= 0;
            conv2d_25_out_page_dma_offset <= 512;
            conv2d_25_out_page <= 0;
          end 
          conv2d_25_prev_row_count <= conv2d_25_row_count;
          conv2d_25_prev_bat_count <= conv2d_25_bat_count;
          conv2d_25_prev_och_count <= conv2d_25_och_count;
          if((conv2d_25_row_count >= cparam_conv2d_25_max_row_count) && (conv2d_25_bat_count >= cparam_conv2d_25_max_bat_count) && (conv2d_25_och_count >= cparam_conv2d_25_max_och_count)) begin
            conv2d_25_skip_read_filter <= 1;
          end 
          if((cparam_conv2d_25_data_stationary == 1) && cparam_conv2d_25_keep_filter) begin
            conv2d_25_skip_read_filter <= 1;
          end 
          if((conv2d_25_row_count >= cparam_conv2d_25_max_row_count) && (conv2d_25_bat_count >= cparam_conv2d_25_max_bat_count) && (conv2d_25_och_count >= cparam_conv2d_25_max_och_count)) begin
            conv2d_25_skip_read_act <= 1;
          end 
          if((cparam_conv2d_25_data_stationary == 0) && (conv2d_25_row_count >= cparam_conv2d_25_max_row_count) && (conv2d_25_bat_count >= cparam_conv2d_25_max_bat_count) && cparam_conv2d_25_keep_input) begin
            conv2d_25_skip_read_act <= 1;
          end 
          if((conv2d_25_row_count >= cparam_conv2d_25_max_row_count) && (conv2d_25_bat_count >= cparam_conv2d_25_max_bat_count) && (conv2d_25_och_count >= cparam_conv2d_25_max_och_count)) begin
            conv2d_25_skip_comp <= 1;
          end 
          if(conv2d_25_skip_write_out && (conv2d_25_prev_row_count == 0) && (conv2d_25_prev_bat_count == 0) && (conv2d_25_prev_och_count == 0)) begin
            conv2d_25_skip_write_out <= 0;
          end 
          if(cparam_conv2d_25_data_stationary == 0) begin
            control_conv2d_25 <= control_conv2d_25_12;
          end 
          if((cparam_conv2d_25_data_stationary == 0) && (conv2d_25_row_count >= cparam_conv2d_25_max_row_count) && (conv2d_25_bat_count >= cparam_conv2d_25_max_bat_count)) begin
            control_conv2d_25 <= control_conv2d_25_7;
          end 
          if(cparam_conv2d_25_data_stationary == 1) begin
            control_conv2d_25 <= control_conv2d_25_7;
          end 
          if((cparam_conv2d_25_data_stationary == 1) && (conv2d_25_och_count >= cparam_conv2d_25_max_och_count)) begin
            control_conv2d_25 <= control_conv2d_25_12;
          end 
          if(!conv2d_25_skip_write_out && (conv2d_25_prev_och_count >= cparam_conv2d_25_max_och_count) && (conv2d_25_prev_row_count >= cparam_conv2d_25_max_row_count) && (conv2d_25_prev_bat_count >= cparam_conv2d_25_max_bat_count)) begin
            control_conv2d_25 <= control_conv2d_25_33;
          end 
        end
        control_conv2d_25_33: begin
          if(_maxi_write_idle && !_maxi_has_outstanding_write) begin
            control_conv2d_25 <= control_conv2d_25_34;
          end 
        end
        control_conv2d_25_34: begin
          if(main_fsm == 14) begin
            _control_conv2d_25_called <= 0;
          end 
          if(main_fsm == 31) begin
            _control_conv2d_25_called <= 0;
          end 
          if(main_fsm == 48) begin
            _control_conv2d_25_called <= 0;
          end 
          if(main_fsm == 65) begin
            _control_conv2d_25_called <= 0;
          end 
          if(main_fsm == 82) begin
            _control_conv2d_25_called <= 0;
          end 
          if(main_fsm == 99) begin
            _control_conv2d_25_called <= 0;
          end 
          if(main_fsm == 115) begin
            _control_conv2d_25_called <= 0;
          end 
          if(main_fsm == 14) begin
            control_conv2d_25 <= control_conv2d_25_init;
          end 
          if(main_fsm == 31) begin
            control_conv2d_25 <= control_conv2d_25_init;
          end 
          if(main_fsm == 48) begin
            control_conv2d_25 <= control_conv2d_25_init;
          end 
          if(main_fsm == 65) begin
            control_conv2d_25 <= control_conv2d_25_init;
          end 
          if(main_fsm == 82) begin
            control_conv2d_25 <= control_conv2d_25_init;
          end 
          if(main_fsm == 99) begin
            control_conv2d_25 <= control_conv2d_25_init;
          end 
          if(main_fsm == 115) begin
            control_conv2d_25 <= control_conv2d_25_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_read_req_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_read_req_fsm <= _maxi_read_req_fsm_init;
      _maxi_read_cont <= 0;
    end else begin
      case(_maxi_read_req_fsm)
        _maxi_read_req_fsm_init: begin
          if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full) begin
            _maxi_read_req_fsm <= _maxi_read_req_fsm_1;
          end 
        end
        _maxi_read_req_fsm_1: begin
          if(maxi_arready || !maxi_arvalid) begin
            _maxi_read_cont <= 1;
          end 
          if((maxi_arready || !maxi_arvalid) && (_maxi_read_global_size == 0)) begin
            _maxi_read_cont <= 0;
          end 
          if(maxi_arready || !maxi_arvalid) begin
            _maxi_read_req_fsm <= _maxi_read_req_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_read_data_fsm_1 = 1;
  localparam _maxi_read_data_fsm_2 = 2;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
    end else begin
      case(_maxi_read_data_fsm)
        _maxi_read_data_fsm_init: begin
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 6)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 7)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 8)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 9)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
        end
        _maxi_read_data_fsm_1: begin
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
        end
        _maxi_read_data_fsm_2: begin
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_0_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_0 <= write_burst_fsm_0_init;
      write_burst_addr_76 <= 0;
      write_burst_stride_77 <= 0;
      write_burst_length_78 <= 0;
      write_burst_done_79 <= 0;
    end else begin
      case(write_burst_fsm_0)
        write_burst_fsm_0_init: begin
          write_burst_addr_76 <= _maxi_read_local_addr_buf;
          write_burst_stride_77 <= _maxi_read_local_stride_buf;
          write_burst_length_78 <= _maxi_read_local_size_buf;
          write_burst_done_79 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 1) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_0 <= write_burst_fsm_0_1;
          end 
        end
        write_burst_fsm_0_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_addr_76 <= write_burst_addr_76 + write_burst_stride_77;
            write_burst_length_78 <= write_burst_length_78 - 1;
            write_burst_done_79 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_78 <= 1)) begin
            write_burst_done_79 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_done_79 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_78 <= 1)) begin
            write_burst_fsm_0 <= write_burst_fsm_0_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_fsm_0 <= write_burst_fsm_0_init;
          end 
          if(0) begin
            write_burst_fsm_0 <= write_burst_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_1_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_1 <= write_burst_fsm_1_init;
      write_burst_addr_82 <= 0;
      write_burst_stride_83 <= 0;
      write_burst_length_84 <= 0;
      write_burst_done_85 <= 0;
    end else begin
      case(write_burst_fsm_1)
        write_burst_fsm_1_init: begin
          write_burst_addr_82 <= _maxi_read_local_addr_buf;
          write_burst_stride_83 <= _maxi_read_local_stride_buf;
          write_burst_length_84 <= _maxi_read_local_size_buf;
          write_burst_done_85 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 2) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_1 <= write_burst_fsm_1_1;
          end 
        end
        write_burst_fsm_1_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_addr_82 <= write_burst_addr_82 + write_burst_stride_83;
            write_burst_length_84 <= write_burst_length_84 - 1;
            write_burst_done_85 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_84 <= 1)) begin
            write_burst_done_85 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_done_85 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_84 <= 1)) begin
            write_burst_fsm_1 <= write_burst_fsm_1_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_fsm_1 <= write_burst_fsm_1_init;
          end 
          if(0) begin
            write_burst_fsm_1 <= write_burst_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_2_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_2 <= write_burst_fsm_2_init;
      write_burst_addr_90 <= 0;
      write_burst_stride_91 <= 0;
      write_burst_length_92 <= 0;
      write_burst_done_93 <= 0;
    end else begin
      case(write_burst_fsm_2)
        write_burst_fsm_2_init: begin
          write_burst_addr_90 <= _maxi_read_local_addr_buf;
          write_burst_stride_91 <= _maxi_read_local_stride_buf;
          write_burst_length_92 <= _maxi_read_local_size_buf;
          write_burst_done_93 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_2 <= write_burst_fsm_2_1;
          end 
        end
        write_burst_fsm_2_1: begin
          if(write_burst_block_ram_wvalid_88) begin
            write_burst_addr_90 <= write_burst_addr_90 + write_burst_stride_91;
            write_burst_length_92 <= write_burst_length_92 - 1;
            write_burst_done_93 <= 0;
          end 
          if(write_burst_block_ram_wvalid_88 && (write_burst_length_92 <= 1)) begin
            write_burst_done_93 <= 1;
          end 
          if(write_burst_block_ram_wvalid_88 && 0) begin
            write_burst_done_93 <= 1;
          end 
          if(write_burst_block_ram_wvalid_88 && (write_burst_length_92 <= 1)) begin
            write_burst_fsm_2 <= write_burst_fsm_2_init;
          end 
          if(write_burst_block_ram_wvalid_88 && 0) begin
            write_burst_fsm_2 <= write_burst_fsm_2_init;
          end 
          if(write_burst_block_ram_wquit_89) begin
            write_burst_fsm_2 <= write_burst_fsm_2_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_3_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_3 <= write_burst_fsm_3_init;
      write_burst_addr_96 <= 0;
      write_burst_stride_97 <= 0;
      write_burst_length_98 <= 0;
      write_burst_done_99 <= 0;
    end else begin
      case(write_burst_fsm_3)
        write_burst_fsm_3_init: begin
          write_burst_addr_96 <= _maxi_read_local_addr_buf;
          write_burst_stride_97 <= _maxi_read_local_stride_buf;
          write_burst_length_98 <= _maxi_read_local_size_buf;
          write_burst_done_99 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_3 <= write_burst_fsm_3_1;
          end 
        end
        write_burst_fsm_3_1: begin
          if(write_burst_block_ram_wvalid_94) begin
            write_burst_addr_96 <= write_burst_addr_96 + write_burst_stride_97;
            write_burst_length_98 <= write_burst_length_98 - 1;
            write_burst_done_99 <= 0;
          end 
          if(write_burst_block_ram_wvalid_94 && (write_burst_length_98 <= 1)) begin
            write_burst_done_99 <= 1;
          end 
          if(write_burst_block_ram_wvalid_94 && 0) begin
            write_burst_done_99 <= 1;
          end 
          if(write_burst_block_ram_wvalid_94 && (write_burst_length_98 <= 1)) begin
            write_burst_fsm_3 <= write_burst_fsm_3_init;
          end 
          if(write_burst_block_ram_wvalid_94 && 0) begin
            write_burst_fsm_3 <= write_burst_fsm_3_init;
          end 
          if(write_burst_block_ram_wquit_95) begin
            write_burst_fsm_3 <= write_burst_fsm_3_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_4_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_4 <= write_burst_fsm_4_init;
      write_burst_addr_102 <= 0;
      write_burst_stride_103 <= 0;
      write_burst_length_104 <= 0;
      write_burst_done_105 <= 0;
    end else begin
      case(write_burst_fsm_4)
        write_burst_fsm_4_init: begin
          write_burst_addr_102 <= _maxi_read_local_addr_buf;
          write_burst_stride_103 <= _maxi_read_local_stride_buf;
          write_burst_length_104 <= _maxi_read_local_size_buf;
          write_burst_done_105 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_4 <= write_burst_fsm_4_1;
          end 
        end
        write_burst_fsm_4_1: begin
          if(write_burst_block_ram_wvalid_100) begin
            write_burst_addr_102 <= write_burst_addr_102 + write_burst_stride_103;
            write_burst_length_104 <= write_burst_length_104 - 1;
            write_burst_done_105 <= 0;
          end 
          if(write_burst_block_ram_wvalid_100 && (write_burst_length_104 <= 1)) begin
            write_burst_done_105 <= 1;
          end 
          if(write_burst_block_ram_wvalid_100 && 0) begin
            write_burst_done_105 <= 1;
          end 
          if(write_burst_block_ram_wvalid_100 && (write_burst_length_104 <= 1)) begin
            write_burst_fsm_4 <= write_burst_fsm_4_init;
          end 
          if(write_burst_block_ram_wvalid_100 && 0) begin
            write_burst_fsm_4 <= write_burst_fsm_4_init;
          end 
          if(write_burst_block_ram_wquit_101) begin
            write_burst_fsm_4 <= write_burst_fsm_4_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_5_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_5 <= write_burst_fsm_5_init;
      write_burst_addr_108 <= 0;
      write_burst_stride_109 <= 0;
      write_burst_length_110 <= 0;
      write_burst_done_111 <= 0;
    end else begin
      case(write_burst_fsm_5)
        write_burst_fsm_5_init: begin
          write_burst_addr_108 <= _maxi_read_local_addr_buf;
          write_burst_stride_109 <= _maxi_read_local_stride_buf;
          write_burst_length_110 <= _maxi_read_local_size_buf;
          write_burst_done_111 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_5 <= write_burst_fsm_5_1;
          end 
        end
        write_burst_fsm_5_1: begin
          if(write_burst_block_ram_wvalid_106) begin
            write_burst_addr_108 <= write_burst_addr_108 + write_burst_stride_109;
            write_burst_length_110 <= write_burst_length_110 - 1;
            write_burst_done_111 <= 0;
          end 
          if(write_burst_block_ram_wvalid_106 && (write_burst_length_110 <= 1)) begin
            write_burst_done_111 <= 1;
          end 
          if(write_burst_block_ram_wvalid_106 && 0) begin
            write_burst_done_111 <= 1;
          end 
          if(write_burst_block_ram_wvalid_106 && (write_burst_length_110 <= 1)) begin
            write_burst_fsm_5 <= write_burst_fsm_5_init;
          end 
          if(write_burst_block_ram_wvalid_106 && 0) begin
            write_burst_fsm_5 <= write_burst_fsm_5_init;
          end 
          if(write_burst_block_ram_wquit_107) begin
            write_burst_fsm_5 <= write_burst_fsm_5_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_6_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_6 <= write_burst_fsm_6_init;
      write_burst_addr_114 <= 0;
      write_burst_stride_115 <= 0;
      write_burst_length_116 <= 0;
      write_burst_done_117 <= 0;
    end else begin
      case(write_burst_fsm_6)
        write_burst_fsm_6_init: begin
          write_burst_addr_114 <= _maxi_read_local_addr_buf;
          write_burst_stride_115 <= _maxi_read_local_stride_buf;
          write_burst_length_116 <= _maxi_read_local_size_buf;
          write_burst_done_117 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_6 <= write_burst_fsm_6_1;
          end 
        end
        write_burst_fsm_6_1: begin
          if(write_burst_block_ram_wvalid_112) begin
            write_burst_addr_114 <= write_burst_addr_114 + write_burst_stride_115;
            write_burst_length_116 <= write_burst_length_116 - 1;
            write_burst_done_117 <= 0;
          end 
          if(write_burst_block_ram_wvalid_112 && (write_burst_length_116 <= 1)) begin
            write_burst_done_117 <= 1;
          end 
          if(write_burst_block_ram_wvalid_112 && 0) begin
            write_burst_done_117 <= 1;
          end 
          if(write_burst_block_ram_wvalid_112 && (write_burst_length_116 <= 1)) begin
            write_burst_fsm_6 <= write_burst_fsm_6_init;
          end 
          if(write_burst_block_ram_wvalid_112 && 0) begin
            write_burst_fsm_6 <= write_burst_fsm_6_init;
          end 
          if(write_burst_block_ram_wquit_113) begin
            write_burst_fsm_6 <= write_burst_fsm_6_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_7_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_7 <= write_burst_fsm_7_init;
      write_burst_addr_120 <= 0;
      write_burst_stride_121 <= 0;
      write_burst_length_122 <= 0;
      write_burst_done_123 <= 0;
    end else begin
      case(write_burst_fsm_7)
        write_burst_fsm_7_init: begin
          write_burst_addr_120 <= _maxi_read_local_addr_buf;
          write_burst_stride_121 <= _maxi_read_local_stride_buf;
          write_burst_length_122 <= _maxi_read_local_size_buf;
          write_burst_done_123 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_7 <= write_burst_fsm_7_1;
          end 
        end
        write_burst_fsm_7_1: begin
          if(write_burst_block_ram_wvalid_118) begin
            write_burst_addr_120 <= write_burst_addr_120 + write_burst_stride_121;
            write_burst_length_122 <= write_burst_length_122 - 1;
            write_burst_done_123 <= 0;
          end 
          if(write_burst_block_ram_wvalid_118 && (write_burst_length_122 <= 1)) begin
            write_burst_done_123 <= 1;
          end 
          if(write_burst_block_ram_wvalid_118 && 0) begin
            write_burst_done_123 <= 1;
          end 
          if(write_burst_block_ram_wvalid_118 && (write_burst_length_122 <= 1)) begin
            write_burst_fsm_7 <= write_burst_fsm_7_init;
          end 
          if(write_burst_block_ram_wvalid_118 && 0) begin
            write_burst_fsm_7 <= write_burst_fsm_7_init;
          end 
          if(write_burst_block_ram_wquit_119) begin
            write_burst_fsm_7 <= write_burst_fsm_7_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_8_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_8 <= write_burst_fsm_8_init;
      write_burst_addr_126 <= 0;
      write_burst_stride_127 <= 0;
      write_burst_length_128 <= 0;
      write_burst_done_129 <= 0;
    end else begin
      case(write_burst_fsm_8)
        write_burst_fsm_8_init: begin
          write_burst_addr_126 <= _maxi_read_local_addr_buf;
          write_burst_stride_127 <= _maxi_read_local_stride_buf;
          write_burst_length_128 <= _maxi_read_local_size_buf;
          write_burst_done_129 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_8 <= write_burst_fsm_8_1;
          end 
        end
        write_burst_fsm_8_1: begin
          if(write_burst_block_ram_wvalid_124) begin
            write_burst_addr_126 <= write_burst_addr_126 + write_burst_stride_127;
            write_burst_length_128 <= write_burst_length_128 - 1;
            write_burst_done_129 <= 0;
          end 
          if(write_burst_block_ram_wvalid_124 && (write_burst_length_128 <= 1)) begin
            write_burst_done_129 <= 1;
          end 
          if(write_burst_block_ram_wvalid_124 && 0) begin
            write_burst_done_129 <= 1;
          end 
          if(write_burst_block_ram_wvalid_124 && (write_burst_length_128 <= 1)) begin
            write_burst_fsm_8 <= write_burst_fsm_8_init;
          end 
          if(write_burst_block_ram_wvalid_124 && 0) begin
            write_burst_fsm_8 <= write_burst_fsm_8_init;
          end 
          if(write_burst_block_ram_wquit_125) begin
            write_burst_fsm_8 <= write_burst_fsm_8_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_9_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_9 <= write_burst_fsm_9_init;
      write_burst_addr_132 <= 0;
      write_burst_stride_133 <= 0;
      write_burst_length_134 <= 0;
      write_burst_done_135 <= 0;
    end else begin
      case(write_burst_fsm_9)
        write_burst_fsm_9_init: begin
          write_burst_addr_132 <= _maxi_read_local_addr_buf;
          write_burst_stride_133 <= _maxi_read_local_stride_buf;
          write_burst_length_134 <= _maxi_read_local_size_buf;
          write_burst_done_135 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_9 <= write_burst_fsm_9_1;
          end 
        end
        write_burst_fsm_9_1: begin
          if(write_burst_block_ram_wvalid_130) begin
            write_burst_addr_132 <= write_burst_addr_132 + write_burst_stride_133;
            write_burst_length_134 <= write_burst_length_134 - 1;
            write_burst_done_135 <= 0;
          end 
          if(write_burst_block_ram_wvalid_130 && (write_burst_length_134 <= 1)) begin
            write_burst_done_135 <= 1;
          end 
          if(write_burst_block_ram_wvalid_130 && 0) begin
            write_burst_done_135 <= 1;
          end 
          if(write_burst_block_ram_wvalid_130 && (write_burst_length_134 <= 1)) begin
            write_burst_fsm_9 <= write_burst_fsm_9_init;
          end 
          if(write_burst_block_ram_wvalid_130 && 0) begin
            write_burst_fsm_9 <= write_burst_fsm_9_init;
          end 
          if(write_burst_block_ram_wquit_131) begin
            write_burst_fsm_9 <= write_burst_fsm_9_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_10_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_10 <= write_burst_fsm_10_init;
      write_burst_addr_138 <= 0;
      write_burst_stride_139 <= 0;
      write_burst_length_140 <= 0;
      write_burst_done_141 <= 0;
    end else begin
      case(write_burst_fsm_10)
        write_burst_fsm_10_init: begin
          write_burst_addr_138 <= _maxi_read_local_addr_buf;
          write_burst_stride_139 <= _maxi_read_local_stride_buf;
          write_burst_length_140 <= _maxi_read_local_size_buf;
          write_burst_done_141 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_10 <= write_burst_fsm_10_1;
          end 
        end
        write_burst_fsm_10_1: begin
          if(write_burst_block_ram_wvalid_136) begin
            write_burst_addr_138 <= write_burst_addr_138 + write_burst_stride_139;
            write_burst_length_140 <= write_burst_length_140 - 1;
            write_burst_done_141 <= 0;
          end 
          if(write_burst_block_ram_wvalid_136 && (write_burst_length_140 <= 1)) begin
            write_burst_done_141 <= 1;
          end 
          if(write_burst_block_ram_wvalid_136 && 0) begin
            write_burst_done_141 <= 1;
          end 
          if(write_burst_block_ram_wvalid_136 && (write_burst_length_140 <= 1)) begin
            write_burst_fsm_10 <= write_burst_fsm_10_init;
          end 
          if(write_burst_block_ram_wvalid_136 && 0) begin
            write_burst_fsm_10 <= write_burst_fsm_10_init;
          end 
          if(write_burst_block_ram_wquit_137) begin
            write_burst_fsm_10 <= write_burst_fsm_10_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_11_1 = 1;
  localparam write_burst_block_fsm_11_2 = 2;
  localparam write_burst_block_fsm_11_3 = 3;
  localparam write_burst_block_fsm_11_4 = 4;
  localparam write_burst_block_fsm_11_5 = 5;
  localparam write_burst_block_fsm_11_6 = 6;
  localparam write_burst_block_fsm_11_7 = 7;
  localparam write_burst_block_fsm_11_8 = 8;
  localparam write_burst_block_fsm_11_9 = 9;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
      write_burst_block_length_142 <= 0;
      write_burst_block_blocksize_143 <= 0;
      write_burst_block_done_144 <= 0;
      write_burst_block_count_145 <= 0;
    end else begin
      case(write_burst_block_fsm_11)
        write_burst_block_fsm_11_init: begin
          write_burst_block_length_142 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_143 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_144 <= 0;
          write_burst_block_count_145 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_1;
          end 
        end
        write_burst_block_fsm_11_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_142 <= write_burst_block_length_142 - 1;
            write_burst_block_done_144 <= 0;
            write_burst_block_count_145 <= write_burst_block_count_145 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_count_145 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_142 <= write_burst_block_length_142 - 1;
            write_burst_block_done_144 <= 0;
            write_burst_block_count_145 <= write_burst_block_count_145 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_count_145 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_142 <= write_burst_block_length_142 - 1;
            write_burst_block_done_144 <= 0;
            write_burst_block_count_145 <= write_burst_block_count_145 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_count_145 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_4;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_4: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_142 <= write_burst_block_length_142 - 1;
            write_burst_block_done_144 <= 0;
            write_burst_block_count_145 <= write_burst_block_count_145 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_count_145 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_5;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_5: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_142 <= write_burst_block_length_142 - 1;
            write_burst_block_done_144 <= 0;
            write_burst_block_count_145 <= write_burst_block_count_145 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_count_145 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_6;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_6: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_142 <= write_burst_block_length_142 - 1;
            write_burst_block_done_144 <= 0;
            write_burst_block_count_145 <= write_burst_block_count_145 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_count_145 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_7;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_7: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_142 <= write_burst_block_length_142 - 1;
            write_burst_block_done_144 <= 0;
            write_burst_block_count_145 <= write_burst_block_count_145 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_count_145 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_8;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_8: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_142 <= write_burst_block_length_142 - 1;
            write_burst_block_done_144 <= 0;
            write_burst_block_count_145 <= write_burst_block_count_145 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_count_145 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_9;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_9: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_142 <= write_burst_block_length_142 - 1;
            write_burst_block_done_144 <= 0;
            write_burst_block_count_145 <= write_burst_block_count_145 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_144 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_count_145 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_145 == write_burst_block_blocksize_143 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_142 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_12_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_12 <= write_burst_fsm_12_init;
      write_burst_addr_150 <= 0;
      write_burst_stride_151 <= 0;
      write_burst_length_152 <= 0;
      write_burst_done_153 <= 0;
    end else begin
      case(write_burst_fsm_12)
        write_burst_fsm_12_init: begin
          write_burst_addr_150 <= _maxi_read_local_addr_buf;
          write_burst_stride_151 <= _maxi_read_local_stride_buf;
          write_burst_length_152 <= _maxi_read_local_size_buf;
          write_burst_done_153 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_12 <= write_burst_fsm_12_1;
          end 
        end
        write_burst_fsm_12_1: begin
          if(write_burst_block_ram_wvalid_148) begin
            write_burst_addr_150 <= write_burst_addr_150 + write_burst_stride_151;
            write_burst_length_152 <= write_burst_length_152 - 1;
            write_burst_done_153 <= 0;
          end 
          if(write_burst_block_ram_wvalid_148 && (write_burst_length_152 <= 1)) begin
            write_burst_done_153 <= 1;
          end 
          if(write_burst_block_ram_wvalid_148 && 0) begin
            write_burst_done_153 <= 1;
          end 
          if(write_burst_block_ram_wvalid_148 && (write_burst_length_152 <= 1)) begin
            write_burst_fsm_12 <= write_burst_fsm_12_init;
          end 
          if(write_burst_block_ram_wvalid_148 && 0) begin
            write_burst_fsm_12 <= write_burst_fsm_12_init;
          end 
          if(write_burst_block_ram_wquit_149) begin
            write_burst_fsm_12 <= write_burst_fsm_12_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_13_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_13 <= write_burst_fsm_13_init;
      write_burst_addr_156 <= 0;
      write_burst_stride_157 <= 0;
      write_burst_length_158 <= 0;
      write_burst_done_159 <= 0;
    end else begin
      case(write_burst_fsm_13)
        write_burst_fsm_13_init: begin
          write_burst_addr_156 <= _maxi_read_local_addr_buf;
          write_burst_stride_157 <= _maxi_read_local_stride_buf;
          write_burst_length_158 <= _maxi_read_local_size_buf;
          write_burst_done_159 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_13 <= write_burst_fsm_13_1;
          end 
        end
        write_burst_fsm_13_1: begin
          if(write_burst_block_ram_wvalid_154) begin
            write_burst_addr_156 <= write_burst_addr_156 + write_burst_stride_157;
            write_burst_length_158 <= write_burst_length_158 - 1;
            write_burst_done_159 <= 0;
          end 
          if(write_burst_block_ram_wvalid_154 && (write_burst_length_158 <= 1)) begin
            write_burst_done_159 <= 1;
          end 
          if(write_burst_block_ram_wvalid_154 && 0) begin
            write_burst_done_159 <= 1;
          end 
          if(write_burst_block_ram_wvalid_154 && (write_burst_length_158 <= 1)) begin
            write_burst_fsm_13 <= write_burst_fsm_13_init;
          end 
          if(write_burst_block_ram_wvalid_154 && 0) begin
            write_burst_fsm_13 <= write_burst_fsm_13_init;
          end 
          if(write_burst_block_ram_wquit_155) begin
            write_burst_fsm_13 <= write_burst_fsm_13_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_14_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_14 <= write_burst_fsm_14_init;
      write_burst_addr_162 <= 0;
      write_burst_stride_163 <= 0;
      write_burst_length_164 <= 0;
      write_burst_done_165 <= 0;
    end else begin
      case(write_burst_fsm_14)
        write_burst_fsm_14_init: begin
          write_burst_addr_162 <= _maxi_read_local_addr_buf;
          write_burst_stride_163 <= _maxi_read_local_stride_buf;
          write_burst_length_164 <= _maxi_read_local_size_buf;
          write_burst_done_165 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_14 <= write_burst_fsm_14_1;
          end 
        end
        write_burst_fsm_14_1: begin
          if(write_burst_block_ram_wvalid_160) begin
            write_burst_addr_162 <= write_burst_addr_162 + write_burst_stride_163;
            write_burst_length_164 <= write_burst_length_164 - 1;
            write_burst_done_165 <= 0;
          end 
          if(write_burst_block_ram_wvalid_160 && (write_burst_length_164 <= 1)) begin
            write_burst_done_165 <= 1;
          end 
          if(write_burst_block_ram_wvalid_160 && 0) begin
            write_burst_done_165 <= 1;
          end 
          if(write_burst_block_ram_wvalid_160 && (write_burst_length_164 <= 1)) begin
            write_burst_fsm_14 <= write_burst_fsm_14_init;
          end 
          if(write_burst_block_ram_wvalid_160 && 0) begin
            write_burst_fsm_14 <= write_burst_fsm_14_init;
          end 
          if(write_burst_block_ram_wquit_161) begin
            write_burst_fsm_14 <= write_burst_fsm_14_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_15_1 = 1;
  localparam write_burst_block_fsm_15_2 = 2;
  localparam write_burst_block_fsm_15_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
      write_burst_block_length_166 <= 0;
      write_burst_block_blocksize_167 <= 0;
      write_burst_block_done_168 <= 0;
      write_burst_block_count_169 <= 0;
    end else begin
      case(write_burst_block_fsm_15)
        write_burst_block_fsm_15_init: begin
          write_burst_block_length_166 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_167 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_168 <= 0;
          write_burst_block_count_169 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_1;
          end 
        end
        write_burst_block_fsm_15_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_166 <= write_burst_block_length_166 - 1;
            write_burst_block_done_168 <= 0;
            write_burst_block_count_169 <= write_burst_block_count_169 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_166 <= 1)) begin
            write_burst_block_done_168 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_168 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_169 == write_burst_block_blocksize_167 - 1)) begin
            write_burst_block_count_169 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_169 == write_burst_block_blocksize_167 - 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_166 <= 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
        end
        write_burst_block_fsm_15_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_166 <= write_burst_block_length_166 - 1;
            write_burst_block_done_168 <= 0;
            write_burst_block_count_169 <= write_burst_block_count_169 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_166 <= 1)) begin
            write_burst_block_done_168 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_168 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_169 == write_burst_block_blocksize_167 - 1)) begin
            write_burst_block_count_169 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_169 == write_burst_block_blocksize_167 - 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_166 <= 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
        end
        write_burst_block_fsm_15_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_166 <= write_burst_block_length_166 - 1;
            write_burst_block_done_168 <= 0;
            write_burst_block_count_169 <= write_burst_block_count_169 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_166 <= 1)) begin
            write_burst_block_done_168 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_168 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_169 == write_burst_block_blocksize_167 - 1)) begin
            write_burst_block_count_169 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_169 == write_burst_block_blocksize_167 - 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_166 <= 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_16_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_16 <= write_burst_fsm_16_init;
      write_burst_addr_174 <= 0;
      write_burst_stride_175 <= 0;
      write_burst_length_176 <= 0;
      write_burst_done_177 <= 0;
    end else begin
      case(write_burst_fsm_16)
        write_burst_fsm_16_init: begin
          write_burst_addr_174 <= _maxi_read_local_addr_buf;
          write_burst_stride_175 <= _maxi_read_local_stride_buf;
          write_burst_length_176 <= _maxi_read_local_size_buf;
          write_burst_done_177 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_16 <= write_burst_fsm_16_1;
          end 
        end
        write_burst_fsm_16_1: begin
          if(write_burst_block_ram_wvalid_172) begin
            write_burst_addr_174 <= write_burst_addr_174 + write_burst_stride_175;
            write_burst_length_176 <= write_burst_length_176 - 1;
            write_burst_done_177 <= 0;
          end 
          if(write_burst_block_ram_wvalid_172 && (write_burst_length_176 <= 1)) begin
            write_burst_done_177 <= 1;
          end 
          if(write_burst_block_ram_wvalid_172 && 0) begin
            write_burst_done_177 <= 1;
          end 
          if(write_burst_block_ram_wvalid_172 && (write_burst_length_176 <= 1)) begin
            write_burst_fsm_16 <= write_burst_fsm_16_init;
          end 
          if(write_burst_block_ram_wvalid_172 && 0) begin
            write_burst_fsm_16 <= write_burst_fsm_16_init;
          end 
          if(write_burst_block_ram_wquit_173) begin
            write_burst_fsm_16 <= write_burst_fsm_16_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_17_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_17 <= write_burst_fsm_17_init;
      write_burst_addr_180 <= 0;
      write_burst_stride_181 <= 0;
      write_burst_length_182 <= 0;
      write_burst_done_183 <= 0;
    end else begin
      case(write_burst_fsm_17)
        write_burst_fsm_17_init: begin
          write_burst_addr_180 <= _maxi_read_local_addr_buf;
          write_burst_stride_181 <= _maxi_read_local_stride_buf;
          write_burst_length_182 <= _maxi_read_local_size_buf;
          write_burst_done_183 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_17 <= write_burst_fsm_17_1;
          end 
        end
        write_burst_fsm_17_1: begin
          if(write_burst_block_ram_wvalid_178) begin
            write_burst_addr_180 <= write_burst_addr_180 + write_burst_stride_181;
            write_burst_length_182 <= write_burst_length_182 - 1;
            write_burst_done_183 <= 0;
          end 
          if(write_burst_block_ram_wvalid_178 && (write_burst_length_182 <= 1)) begin
            write_burst_done_183 <= 1;
          end 
          if(write_burst_block_ram_wvalid_178 && 0) begin
            write_burst_done_183 <= 1;
          end 
          if(write_burst_block_ram_wvalid_178 && (write_burst_length_182 <= 1)) begin
            write_burst_fsm_17 <= write_burst_fsm_17_init;
          end 
          if(write_burst_block_ram_wvalid_178 && 0) begin
            write_burst_fsm_17 <= write_burst_fsm_17_init;
          end 
          if(write_burst_block_ram_wquit_179) begin
            write_burst_fsm_17 <= write_burst_fsm_17_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_18_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_18 <= write_burst_fsm_18_init;
      write_burst_addr_186 <= 0;
      write_burst_stride_187 <= 0;
      write_burst_length_188 <= 0;
      write_burst_done_189 <= 0;
    end else begin
      case(write_burst_fsm_18)
        write_burst_fsm_18_init: begin
          write_burst_addr_186 <= _maxi_read_local_addr_buf;
          write_burst_stride_187 <= _maxi_read_local_stride_buf;
          write_burst_length_188 <= _maxi_read_local_size_buf;
          write_burst_done_189 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_18 <= write_burst_fsm_18_1;
          end 
        end
        write_burst_fsm_18_1: begin
          if(write_burst_block_ram_wvalid_184) begin
            write_burst_addr_186 <= write_burst_addr_186 + write_burst_stride_187;
            write_burst_length_188 <= write_burst_length_188 - 1;
            write_burst_done_189 <= 0;
          end 
          if(write_burst_block_ram_wvalid_184 && (write_burst_length_188 <= 1)) begin
            write_burst_done_189 <= 1;
          end 
          if(write_burst_block_ram_wvalid_184 && 0) begin
            write_burst_done_189 <= 1;
          end 
          if(write_burst_block_ram_wvalid_184 && (write_burst_length_188 <= 1)) begin
            write_burst_fsm_18 <= write_burst_fsm_18_init;
          end 
          if(write_burst_block_ram_wvalid_184 && 0) begin
            write_burst_fsm_18 <= write_burst_fsm_18_init;
          end 
          if(write_burst_block_ram_wquit_185) begin
            write_burst_fsm_18 <= write_burst_fsm_18_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_19_1 = 1;
  localparam write_burst_block_fsm_19_2 = 2;
  localparam write_burst_block_fsm_19_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
      write_burst_block_length_190 <= 0;
      write_burst_block_blocksize_191 <= 0;
      write_burst_block_done_192 <= 0;
      write_burst_block_count_193 <= 0;
    end else begin
      case(write_burst_block_fsm_19)
        write_burst_block_fsm_19_init: begin
          write_burst_block_length_190 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_191 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_192 <= 0;
          write_burst_block_count_193 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_1;
          end 
        end
        write_burst_block_fsm_19_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_190 <= write_burst_block_length_190 - 1;
            write_burst_block_done_192 <= 0;
            write_burst_block_count_193 <= write_burst_block_count_193 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_190 <= 1)) begin
            write_burst_block_done_192 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_192 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_193 == write_burst_block_blocksize_191 - 1)) begin
            write_burst_block_count_193 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_193 == write_burst_block_blocksize_191 - 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_190 <= 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
        end
        write_burst_block_fsm_19_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_190 <= write_burst_block_length_190 - 1;
            write_burst_block_done_192 <= 0;
            write_burst_block_count_193 <= write_burst_block_count_193 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_190 <= 1)) begin
            write_burst_block_done_192 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_192 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_193 == write_burst_block_blocksize_191 - 1)) begin
            write_burst_block_count_193 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_193 == write_burst_block_blocksize_191 - 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_190 <= 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
        end
        write_burst_block_fsm_19_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_190 <= write_burst_block_length_190 - 1;
            write_burst_block_done_192 <= 0;
            write_burst_block_count_193 <= write_burst_block_count_193 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_190 <= 1)) begin
            write_burst_block_done_192 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_192 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_193 == write_burst_block_blocksize_191 - 1)) begin
            write_burst_block_count_193 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_193 == write_burst_block_blocksize_191 - 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_190 <= 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_20_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_20 <= write_burst_fsm_20_init;
      write_burst_addr_198 <= 0;
      write_burst_stride_199 <= 0;
      write_burst_length_200 <= 0;
      write_burst_done_201 <= 0;
    end else begin
      case(write_burst_fsm_20)
        write_burst_fsm_20_init: begin
          write_burst_addr_198 <= _maxi_read_local_addr_buf;
          write_burst_stride_199 <= _maxi_read_local_stride_buf;
          write_burst_length_200 <= _maxi_read_local_size_buf;
          write_burst_done_201 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_20 <= write_burst_fsm_20_1;
          end 
        end
        write_burst_fsm_20_1: begin
          if(write_burst_block_ram_wvalid_196) begin
            write_burst_addr_198 <= write_burst_addr_198 + write_burst_stride_199;
            write_burst_length_200 <= write_burst_length_200 - 1;
            write_burst_done_201 <= 0;
          end 
          if(write_burst_block_ram_wvalid_196 && (write_burst_length_200 <= 1)) begin
            write_burst_done_201 <= 1;
          end 
          if(write_burst_block_ram_wvalid_196 && 0) begin
            write_burst_done_201 <= 1;
          end 
          if(write_burst_block_ram_wvalid_196 && (write_burst_length_200 <= 1)) begin
            write_burst_fsm_20 <= write_burst_fsm_20_init;
          end 
          if(write_burst_block_ram_wvalid_196 && 0) begin
            write_burst_fsm_20 <= write_burst_fsm_20_init;
          end 
          if(write_burst_block_ram_wquit_197) begin
            write_burst_fsm_20 <= write_burst_fsm_20_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_21_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_21 <= write_burst_fsm_21_init;
      write_burst_addr_204 <= 0;
      write_burst_stride_205 <= 0;
      write_burst_length_206 <= 0;
      write_burst_done_207 <= 0;
    end else begin
      case(write_burst_fsm_21)
        write_burst_fsm_21_init: begin
          write_burst_addr_204 <= _maxi_read_local_addr_buf;
          write_burst_stride_205 <= _maxi_read_local_stride_buf;
          write_burst_length_206 <= _maxi_read_local_size_buf;
          write_burst_done_207 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_21 <= write_burst_fsm_21_1;
          end 
        end
        write_burst_fsm_21_1: begin
          if(write_burst_block_ram_wvalid_202) begin
            write_burst_addr_204 <= write_burst_addr_204 + write_burst_stride_205;
            write_burst_length_206 <= write_burst_length_206 - 1;
            write_burst_done_207 <= 0;
          end 
          if(write_burst_block_ram_wvalid_202 && (write_burst_length_206 <= 1)) begin
            write_burst_done_207 <= 1;
          end 
          if(write_burst_block_ram_wvalid_202 && 0) begin
            write_burst_done_207 <= 1;
          end 
          if(write_burst_block_ram_wvalid_202 && (write_burst_length_206 <= 1)) begin
            write_burst_fsm_21 <= write_burst_fsm_21_init;
          end 
          if(write_burst_block_ram_wvalid_202 && 0) begin
            write_burst_fsm_21 <= write_burst_fsm_21_init;
          end 
          if(write_burst_block_ram_wquit_203) begin
            write_burst_fsm_21 <= write_burst_fsm_21_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_22_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_22 <= write_burst_fsm_22_init;
      write_burst_addr_210 <= 0;
      write_burst_stride_211 <= 0;
      write_burst_length_212 <= 0;
      write_burst_done_213 <= 0;
    end else begin
      case(write_burst_fsm_22)
        write_burst_fsm_22_init: begin
          write_burst_addr_210 <= _maxi_read_local_addr_buf;
          write_burst_stride_211 <= _maxi_read_local_stride_buf;
          write_burst_length_212 <= _maxi_read_local_size_buf;
          write_burst_done_213 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_22 <= write_burst_fsm_22_1;
          end 
        end
        write_burst_fsm_22_1: begin
          if(write_burst_block_ram_wvalid_208) begin
            write_burst_addr_210 <= write_burst_addr_210 + write_burst_stride_211;
            write_burst_length_212 <= write_burst_length_212 - 1;
            write_burst_done_213 <= 0;
          end 
          if(write_burst_block_ram_wvalid_208 && (write_burst_length_212 <= 1)) begin
            write_burst_done_213 <= 1;
          end 
          if(write_burst_block_ram_wvalid_208 && 0) begin
            write_burst_done_213 <= 1;
          end 
          if(write_burst_block_ram_wvalid_208 && (write_burst_length_212 <= 1)) begin
            write_burst_fsm_22 <= write_burst_fsm_22_init;
          end 
          if(write_burst_block_ram_wvalid_208 && 0) begin
            write_burst_fsm_22 <= write_burst_fsm_22_init;
          end 
          if(write_burst_block_ram_wquit_209) begin
            write_burst_fsm_22 <= write_burst_fsm_22_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_23_1 = 1;
  localparam write_burst_block_fsm_23_2 = 2;
  localparam write_burst_block_fsm_23_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
      write_burst_block_length_214 <= 0;
      write_burst_block_blocksize_215 <= 0;
      write_burst_block_done_216 <= 0;
      write_burst_block_count_217 <= 0;
    end else begin
      case(write_burst_block_fsm_23)
        write_burst_block_fsm_23_init: begin
          write_burst_block_length_214 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_215 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_216 <= 0;
          write_burst_block_count_217 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_1;
          end 
        end
        write_burst_block_fsm_23_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_214 <= write_burst_block_length_214 - 1;
            write_burst_block_done_216 <= 0;
            write_burst_block_count_217 <= write_burst_block_count_217 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_214 <= 1)) begin
            write_burst_block_done_216 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_216 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_217 == write_burst_block_blocksize_215 - 1)) begin
            write_burst_block_count_217 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_217 == write_burst_block_blocksize_215 - 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_214 <= 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
        end
        write_burst_block_fsm_23_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_214 <= write_burst_block_length_214 - 1;
            write_burst_block_done_216 <= 0;
            write_burst_block_count_217 <= write_burst_block_count_217 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_214 <= 1)) begin
            write_burst_block_done_216 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_216 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_217 == write_burst_block_blocksize_215 - 1)) begin
            write_burst_block_count_217 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_217 == write_burst_block_blocksize_215 - 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_214 <= 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
        end
        write_burst_block_fsm_23_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_214 <= write_burst_block_length_214 - 1;
            write_burst_block_done_216 <= 0;
            write_burst_block_count_217 <= write_burst_block_count_217 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_214 <= 1)) begin
            write_burst_block_done_216 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_216 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_217 == write_burst_block_blocksize_215 - 1)) begin
            write_burst_block_count_217 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_217 == write_burst_block_blocksize_215 - 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_214 <= 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
        end
      endcase
    end
  end

  localparam conv2d_25_comp_fsm_1 = 1;
  localparam conv2d_25_comp_fsm_2 = 2;
  localparam conv2d_25_comp_fsm_3 = 3;
  localparam conv2d_25_comp_fsm_4 = 4;
  localparam conv2d_25_comp_fsm_5 = 5;
  localparam conv2d_25_comp_fsm_6 = 6;

  always @(posedge CLK) begin
    if(RST) begin
      conv2d_25_comp_fsm <= conv2d_25_comp_fsm_init;
      conv2d_25_stream_act_local_0 <= 0;
      conv2d_25_stream_act_local_1 <= 0;
      conv2d_25_stream_act_local_2 <= 0;
      conv2d_25_stream_act_local_3 <= 0;
      conv2d_25_stream_act_local_4 <= 0;
      conv2d_25_stream_act_local_5 <= 0;
      conv2d_25_stream_act_local_6 <= 0;
      conv2d_25_stream_act_local_7 <= 0;
      conv2d_25_stream_act_local_8 <= 0;
      conv2d_25_stream_out_local_col <= 0;
      conv2d_25_stream_out_local_val <= 0;
      conv2d_25_col_count <= 0;
      conv2d_25_col_select <= 0;
      conv2d_25_filter_page_comp_offset_buf <= 0;
      conv2d_25_act_page_comp_offset_buf_0 <= 0;
      conv2d_25_act_page_comp_offset_buf_1 <= 0;
      conv2d_25_act_page_comp_offset_buf_2 <= 0;
      conv2d_25_out_page_comp_offset_buf <= 0;
      conv2d_25_row_count_buf <= 0;
      conv2d_25_row_select_buf <= 0;
      conv2d_25_och_count_buf <= 0;
      conv2d_25_next_stream_num_ops <= 0;
      conv2d_25_stream_pad_masks <= 0;
      conv2d_25_sync_comp_count <= 0;
    end else begin
      if(_stream_conv2d_25_sink_stop) begin
        conv2d_25_sync_comp_count <= conv2d_25_sync_comp_count + 1;
      end 
      if(control_conv2d_25 == 6) begin
        conv2d_25_sync_comp_count <= 0;
      end 
      case(conv2d_25_comp_fsm)
        conv2d_25_comp_fsm_init: begin
          if((control_conv2d_25 == 25) && !conv2d_25_skip_comp) begin
            conv2d_25_comp_fsm <= conv2d_25_comp_fsm_1;
          end 
        end
        conv2d_25_comp_fsm_1: begin
          conv2d_25_stream_act_local_0 <= 0;
          if(cparam_conv2d_25_stream_act_local_small_flags_0) begin
            conv2d_25_stream_act_local_0 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_25_stream_act_local_large_flags_0) begin
            conv2d_25_stream_act_local_0 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          conv2d_25_stream_act_local_1 <= 0;
          if(cparam_conv2d_25_stream_act_local_small_flags_1) begin
            conv2d_25_stream_act_local_1 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_25_stream_act_local_large_flags_1) begin
            conv2d_25_stream_act_local_1 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          conv2d_25_stream_act_local_2 <= 0;
          if(cparam_conv2d_25_stream_act_local_small_flags_2) begin
            conv2d_25_stream_act_local_2 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_25_stream_act_local_large_flags_2) begin
            conv2d_25_stream_act_local_2 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          conv2d_25_stream_act_local_3 <= 0;
          if(cparam_conv2d_25_stream_act_local_small_flags_0) begin
            conv2d_25_stream_act_local_3 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_25_stream_act_local_large_flags_0) begin
            conv2d_25_stream_act_local_3 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          conv2d_25_stream_act_local_4 <= 0;
          if(cparam_conv2d_25_stream_act_local_small_flags_1) begin
            conv2d_25_stream_act_local_4 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_25_stream_act_local_large_flags_1) begin
            conv2d_25_stream_act_local_4 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          conv2d_25_stream_act_local_5 <= 0;
          if(cparam_conv2d_25_stream_act_local_small_flags_2) begin
            conv2d_25_stream_act_local_5 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_25_stream_act_local_large_flags_2) begin
            conv2d_25_stream_act_local_5 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          conv2d_25_stream_act_local_6 <= 0;
          if(cparam_conv2d_25_stream_act_local_small_flags_0) begin
            conv2d_25_stream_act_local_6 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_25_stream_act_local_large_flags_0) begin
            conv2d_25_stream_act_local_6 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          conv2d_25_stream_act_local_7 <= 0;
          if(cparam_conv2d_25_stream_act_local_small_flags_1) begin
            conv2d_25_stream_act_local_7 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_25_stream_act_local_large_flags_1) begin
            conv2d_25_stream_act_local_7 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          conv2d_25_stream_act_local_8 <= 0;
          if(cparam_conv2d_25_stream_act_local_small_flags_2) begin
            conv2d_25_stream_act_local_8 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_25_stream_act_local_large_flags_2) begin
            conv2d_25_stream_act_local_8 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          conv2d_25_stream_out_local_col <= 0;
          if((cparam_conv2d_25_data_stationary == 1) && (conv2d_25_och_count == 0)) begin
            conv2d_25_stream_out_local_val <= 0;
          end 
          conv2d_25_col_count <= 0;
          conv2d_25_col_select <= cparam_conv2d_25_col_select_initval;
          conv2d_25_filter_page_comp_offset_buf <= conv2d_25_filter_page_comp_offset;
          conv2d_25_act_page_comp_offset_buf_0 <= conv2d_25_act_page_comp_offset_0;
          conv2d_25_act_page_comp_offset_buf_1 <= conv2d_25_act_page_comp_offset_1;
          conv2d_25_act_page_comp_offset_buf_2 <= conv2d_25_act_page_comp_offset_2;
          conv2d_25_out_page_comp_offset_buf <= conv2d_25_out_page_comp_offset;
          conv2d_25_row_count_buf <= conv2d_25_row_count;
          conv2d_25_row_select_buf <= conv2d_25_row_select;
          conv2d_25_och_count_buf <= conv2d_25_och_count;
          conv2d_25_next_stream_num_ops <= (conv2d_25_och_count >= cparam_conv2d_25_max_och_count)? cparam_conv2d_25_stream_num_ops_res : cparam_conv2d_25_stream_num_ops;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_2;
        end
        conv2d_25_comp_fsm_2: begin
          conv2d_25_stream_pad_masks <= { conv2d_25_stream_pad_mask_2_2, conv2d_25_stream_pad_mask_2_1, conv2d_25_stream_pad_mask_2_0, conv2d_25_stream_pad_mask_1_2, conv2d_25_stream_pad_mask_1_1, conv2d_25_stream_pad_mask_1_0, conv2d_25_stream_pad_mask_0_2, conv2d_25_stream_pad_mask_0_1, conv2d_25_stream_pad_mask_0_0 };
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_3;
        end
        conv2d_25_comp_fsm_3: begin
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          if(_stream_conv2d_25_stream_oready) begin
            conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
          end 
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_4;
        end
        conv2d_25_comp_fsm_4: begin
          if(!_stream_conv2d_25_source_busy) begin
            conv2d_25_comp_fsm <= conv2d_25_comp_fsm_5;
          end 
        end
        conv2d_25_comp_fsm_5: begin
          if(_stream_conv2d_25_busy) begin
            conv2d_25_comp_fsm <= conv2d_25_comp_fsm_6;
          end 
        end
        conv2d_25_comp_fsm_6: begin
          if(!((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_0 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_1 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_2 : 0)) begin
            conv2d_25_stream_act_local_0 <= conv2d_25_stream_act_local_0 + cparam_conv2d_25_inc_act_laddr_small;
          end 
          if((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_0 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_1 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_2 : 0) begin
            conv2d_25_stream_act_local_0 <= conv2d_25_stream_act_local_0 + cparam_conv2d_25_inc_act_laddr_large;
          end 
          if(conv2d_25_col_count >= cparam_conv2d_25_max_col_count) begin
            conv2d_25_stream_act_local_0 <= 0;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_small_flags_0) begin
            conv2d_25_stream_act_local_0 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_large_flags_0) begin
            conv2d_25_stream_act_local_0 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          if(!((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_3 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_4 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_5 : 0)) begin
            conv2d_25_stream_act_local_1 <= conv2d_25_stream_act_local_1 + cparam_conv2d_25_inc_act_laddr_small;
          end 
          if((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_3 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_4 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_5 : 0) begin
            conv2d_25_stream_act_local_1 <= conv2d_25_stream_act_local_1 + cparam_conv2d_25_inc_act_laddr_large;
          end 
          if(conv2d_25_col_count >= cparam_conv2d_25_max_col_count) begin
            conv2d_25_stream_act_local_1 <= 0;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_small_flags_1) begin
            conv2d_25_stream_act_local_1 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_large_flags_1) begin
            conv2d_25_stream_act_local_1 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          if(!((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_6 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_7 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_8 : 0)) begin
            conv2d_25_stream_act_local_2 <= conv2d_25_stream_act_local_2 + cparam_conv2d_25_inc_act_laddr_small;
          end 
          if((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_6 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_7 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_8 : 0) begin
            conv2d_25_stream_act_local_2 <= conv2d_25_stream_act_local_2 + cparam_conv2d_25_inc_act_laddr_large;
          end 
          if(conv2d_25_col_count >= cparam_conv2d_25_max_col_count) begin
            conv2d_25_stream_act_local_2 <= 0;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_small_flags_2) begin
            conv2d_25_stream_act_local_2 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_large_flags_2) begin
            conv2d_25_stream_act_local_2 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          if(!((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_9 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_10 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_11 : 0)) begin
            conv2d_25_stream_act_local_3 <= conv2d_25_stream_act_local_3 + cparam_conv2d_25_inc_act_laddr_small;
          end 
          if((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_9 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_10 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_11 : 0) begin
            conv2d_25_stream_act_local_3 <= conv2d_25_stream_act_local_3 + cparam_conv2d_25_inc_act_laddr_large;
          end 
          if(conv2d_25_col_count >= cparam_conv2d_25_max_col_count) begin
            conv2d_25_stream_act_local_3 <= 0;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_small_flags_0) begin
            conv2d_25_stream_act_local_3 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_large_flags_0) begin
            conv2d_25_stream_act_local_3 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          if(!((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_12 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_13 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_14 : 0)) begin
            conv2d_25_stream_act_local_4 <= conv2d_25_stream_act_local_4 + cparam_conv2d_25_inc_act_laddr_small;
          end 
          if((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_12 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_13 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_14 : 0) begin
            conv2d_25_stream_act_local_4 <= conv2d_25_stream_act_local_4 + cparam_conv2d_25_inc_act_laddr_large;
          end 
          if(conv2d_25_col_count >= cparam_conv2d_25_max_col_count) begin
            conv2d_25_stream_act_local_4 <= 0;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_small_flags_1) begin
            conv2d_25_stream_act_local_4 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_large_flags_1) begin
            conv2d_25_stream_act_local_4 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          if(!((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_15 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_16 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_17 : 0)) begin
            conv2d_25_stream_act_local_5 <= conv2d_25_stream_act_local_5 + cparam_conv2d_25_inc_act_laddr_small;
          end 
          if((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_15 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_16 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_17 : 0) begin
            conv2d_25_stream_act_local_5 <= conv2d_25_stream_act_local_5 + cparam_conv2d_25_inc_act_laddr_large;
          end 
          if(conv2d_25_col_count >= cparam_conv2d_25_max_col_count) begin
            conv2d_25_stream_act_local_5 <= 0;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_small_flags_2) begin
            conv2d_25_stream_act_local_5 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_large_flags_2) begin
            conv2d_25_stream_act_local_5 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          if(!((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_18 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_19 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_20 : 0)) begin
            conv2d_25_stream_act_local_6 <= conv2d_25_stream_act_local_6 + cparam_conv2d_25_inc_act_laddr_small;
          end 
          if((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_18 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_19 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_20 : 0) begin
            conv2d_25_stream_act_local_6 <= conv2d_25_stream_act_local_6 + cparam_conv2d_25_inc_act_laddr_large;
          end 
          if(conv2d_25_col_count >= cparam_conv2d_25_max_col_count) begin
            conv2d_25_stream_act_local_6 <= 0;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_small_flags_0) begin
            conv2d_25_stream_act_local_6 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_large_flags_0) begin
            conv2d_25_stream_act_local_6 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          if(!((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_21 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_22 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_23 : 0)) begin
            conv2d_25_stream_act_local_7 <= conv2d_25_stream_act_local_7 + cparam_conv2d_25_inc_act_laddr_small;
          end 
          if((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_21 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_22 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_23 : 0) begin
            conv2d_25_stream_act_local_7 <= conv2d_25_stream_act_local_7 + cparam_conv2d_25_inc_act_laddr_large;
          end 
          if(conv2d_25_col_count >= cparam_conv2d_25_max_col_count) begin
            conv2d_25_stream_act_local_7 <= 0;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_small_flags_1) begin
            conv2d_25_stream_act_local_7 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_large_flags_1) begin
            conv2d_25_stream_act_local_7 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          if(!((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_24 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_25 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_26 : 0)) begin
            conv2d_25_stream_act_local_8 <= conv2d_25_stream_act_local_8 + cparam_conv2d_25_inc_act_laddr_small;
          end 
          if((conv2d_25_col_select == 0)? cparam_conv2d_25_inc_act_laddr_conds_24 : 
          (conv2d_25_col_select == 1)? cparam_conv2d_25_inc_act_laddr_conds_25 : 
          (conv2d_25_col_select == 2)? cparam_conv2d_25_inc_act_laddr_conds_26 : 0) begin
            conv2d_25_stream_act_local_8 <= conv2d_25_stream_act_local_8 + cparam_conv2d_25_inc_act_laddr_large;
          end 
          if(conv2d_25_col_count >= cparam_conv2d_25_max_col_count) begin
            conv2d_25_stream_act_local_8 <= 0;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_small_flags_2) begin
            conv2d_25_stream_act_local_8 <= cparam_conv2d_25_stream_act_local_small_offset;
          end 
          if((conv2d_25_col_count >= cparam_conv2d_25_max_col_count) && cparam_conv2d_25_stream_act_local_large_flags_2) begin
            conv2d_25_stream_act_local_8 <= cparam_conv2d_25_stream_act_local_large_offset;
          end 
          if(cparam_conv2d_25_data_stationary == 0) begin
            conv2d_25_stream_out_local_col <= conv2d_25_stream_out_local_col + conv2d_25_next_stream_num_ops;
          end 
          if((cparam_conv2d_25_data_stationary == 0) && (conv2d_25_col_count >= cparam_conv2d_25_max_col_count)) begin
            conv2d_25_stream_out_local_col <= 0;
          end 
          if(cparam_conv2d_25_data_stationary == 1) begin
            conv2d_25_stream_out_local_col <= conv2d_25_stream_out_local_col + cparam_conv2d_25_inc_out_laddr_col;
          end 
          if((cparam_conv2d_25_data_stationary == 1) && (conv2d_25_col_count >= cparam_conv2d_25_max_col_count)) begin
            conv2d_25_stream_out_local_val <= conv2d_25_stream_out_local_val + conv2d_25_next_stream_num_ops;
            conv2d_25_stream_out_local_col <= 0;
          end 
          conv2d_25_col_count <= conv2d_25_col_count + cparam_conv2d_25_stride_col_par_col;
          if(conv2d_25_col_count >= cparam_conv2d_25_max_col_count) begin
            conv2d_25_col_count <= 0;
          end 
          conv2d_25_col_select <= conv2d_25_col_select + cparam_conv2d_25_stride_col_mod_filter_num;
          if(conv2d_25_col_select + cparam_conv2d_25_stride_col_mod_filter_num >= 3) begin
            conv2d_25_col_select <= conv2d_25_col_select - cparam_conv2d_25_filter_num_col_minus_stride_col_mod;
          end 
          if(conv2d_25_col_count >= cparam_conv2d_25_max_col_count) begin
            conv2d_25_col_select <= cparam_conv2d_25_col_select_initval;
          end 
          conv2d_25_comp_fsm <= conv2d_25_comp_fsm_2;
          if(conv2d_25_col_count >= cparam_conv2d_25_max_col_count) begin
            conv2d_25_comp_fsm <= conv2d_25_comp_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_7_source_pat_fsm_0_1 = 1;
  localparam _stream_conv2d_25_source_7_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_7_source_pat_fsm_0 <= _stream_conv2d_25_source_7_source_pat_fsm_0_init;
    end else begin
      case(_stream_conv2d_25_source_7_source_pat_fsm_0)
        _stream_conv2d_25_source_7_source_pat_fsm_0_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_7_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_7_source_pat_fsm_0 <= _stream_conv2d_25_source_7_source_pat_fsm_0_1;
          end 
        end
        _stream_conv2d_25_source_7_source_pat_fsm_0_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_7_source_pat_fsm_0 <= _stream_conv2d_25_source_7_source_pat_fsm_0_init;
          end 
          if((_source_stream_conv2d_25_source_7_pat_count_0 == 0) && (_source_stream_conv2d_25_source_7_pat_count_1 == 0) && (_source_stream_conv2d_25_source_7_pat_count_2 == 0) && (_source_stream_conv2d_25_source_7_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_7_source_pat_fsm_0 <= _stream_conv2d_25_source_7_source_pat_fsm_0_2;
          end 
        end
        _stream_conv2d_25_source_7_source_pat_fsm_0_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_7_source_pat_fsm_0 <= _stream_conv2d_25_source_7_source_pat_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_9_source_pat_fsm_1_1 = 1;
  localparam _stream_conv2d_25_source_9_source_pat_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_9_source_pat_fsm_1 <= _stream_conv2d_25_source_9_source_pat_fsm_1_init;
    end else begin
      case(_stream_conv2d_25_source_9_source_pat_fsm_1)
        _stream_conv2d_25_source_9_source_pat_fsm_1_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_9_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_9_source_pat_fsm_1 <= _stream_conv2d_25_source_9_source_pat_fsm_1_1;
          end 
        end
        _stream_conv2d_25_source_9_source_pat_fsm_1_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_9_source_pat_fsm_1 <= _stream_conv2d_25_source_9_source_pat_fsm_1_init;
          end 
          if((_source_stream_conv2d_25_source_9_pat_count_0 == 0) && (_source_stream_conv2d_25_source_9_pat_count_1 == 0) && (_source_stream_conv2d_25_source_9_pat_count_2 == 0) && (_source_stream_conv2d_25_source_9_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_9_source_pat_fsm_1 <= _stream_conv2d_25_source_9_source_pat_fsm_1_2;
          end 
        end
        _stream_conv2d_25_source_9_source_pat_fsm_1_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_9_source_pat_fsm_1 <= _stream_conv2d_25_source_9_source_pat_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_20_source_pat_fsm_2_1 = 1;
  localparam _stream_conv2d_25_source_20_source_pat_fsm_2_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_20_source_pat_fsm_2 <= _stream_conv2d_25_source_20_source_pat_fsm_2_init;
    end else begin
      case(_stream_conv2d_25_source_20_source_pat_fsm_2)
        _stream_conv2d_25_source_20_source_pat_fsm_2_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_20_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_20_source_pat_fsm_2 <= _stream_conv2d_25_source_20_source_pat_fsm_2_1;
          end 
        end
        _stream_conv2d_25_source_20_source_pat_fsm_2_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_20_source_pat_fsm_2 <= _stream_conv2d_25_source_20_source_pat_fsm_2_init;
          end 
          if((_source_stream_conv2d_25_source_20_pat_count_0 == 0) && (_source_stream_conv2d_25_source_20_pat_count_1 == 0) && (_source_stream_conv2d_25_source_20_pat_count_2 == 0) && (_source_stream_conv2d_25_source_20_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_20_source_pat_fsm_2 <= _stream_conv2d_25_source_20_source_pat_fsm_2_2;
          end 
        end
        _stream_conv2d_25_source_20_source_pat_fsm_2_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_20_source_pat_fsm_2 <= _stream_conv2d_25_source_20_source_pat_fsm_2_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_21_source_pat_fsm_3_1 = 1;
  localparam _stream_conv2d_25_source_21_source_pat_fsm_3_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_21_source_pat_fsm_3 <= _stream_conv2d_25_source_21_source_pat_fsm_3_init;
    end else begin
      case(_stream_conv2d_25_source_21_source_pat_fsm_3)
        _stream_conv2d_25_source_21_source_pat_fsm_3_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_21_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_21_source_pat_fsm_3 <= _stream_conv2d_25_source_21_source_pat_fsm_3_1;
          end 
        end
        _stream_conv2d_25_source_21_source_pat_fsm_3_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_21_source_pat_fsm_3 <= _stream_conv2d_25_source_21_source_pat_fsm_3_init;
          end 
          if((_source_stream_conv2d_25_source_21_pat_count_0 == 0) && (_source_stream_conv2d_25_source_21_pat_count_1 == 0) && (_source_stream_conv2d_25_source_21_pat_count_2 == 0) && (_source_stream_conv2d_25_source_21_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_21_source_pat_fsm_3 <= _stream_conv2d_25_source_21_source_pat_fsm_3_2;
          end 
        end
        _stream_conv2d_25_source_21_source_pat_fsm_3_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_21_source_pat_fsm_3 <= _stream_conv2d_25_source_21_source_pat_fsm_3_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_22_source_pat_fsm_4_1 = 1;
  localparam _stream_conv2d_25_source_22_source_pat_fsm_4_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_22_source_pat_fsm_4 <= _stream_conv2d_25_source_22_source_pat_fsm_4_init;
    end else begin
      case(_stream_conv2d_25_source_22_source_pat_fsm_4)
        _stream_conv2d_25_source_22_source_pat_fsm_4_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_22_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_22_source_pat_fsm_4 <= _stream_conv2d_25_source_22_source_pat_fsm_4_1;
          end 
        end
        _stream_conv2d_25_source_22_source_pat_fsm_4_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_22_source_pat_fsm_4 <= _stream_conv2d_25_source_22_source_pat_fsm_4_init;
          end 
          if((_source_stream_conv2d_25_source_22_pat_count_0 == 0) && (_source_stream_conv2d_25_source_22_pat_count_1 == 0) && (_source_stream_conv2d_25_source_22_pat_count_2 == 0) && (_source_stream_conv2d_25_source_22_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_22_source_pat_fsm_4 <= _stream_conv2d_25_source_22_source_pat_fsm_4_2;
          end 
        end
        _stream_conv2d_25_source_22_source_pat_fsm_4_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_22_source_pat_fsm_4 <= _stream_conv2d_25_source_22_source_pat_fsm_4_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_23_source_pat_fsm_5_1 = 1;
  localparam _stream_conv2d_25_source_23_source_pat_fsm_5_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_23_source_pat_fsm_5 <= _stream_conv2d_25_source_23_source_pat_fsm_5_init;
    end else begin
      case(_stream_conv2d_25_source_23_source_pat_fsm_5)
        _stream_conv2d_25_source_23_source_pat_fsm_5_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_23_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_23_source_pat_fsm_5 <= _stream_conv2d_25_source_23_source_pat_fsm_5_1;
          end 
        end
        _stream_conv2d_25_source_23_source_pat_fsm_5_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_23_source_pat_fsm_5 <= _stream_conv2d_25_source_23_source_pat_fsm_5_init;
          end 
          if((_source_stream_conv2d_25_source_23_pat_count_0 == 0) && (_source_stream_conv2d_25_source_23_pat_count_1 == 0) && (_source_stream_conv2d_25_source_23_pat_count_2 == 0) && (_source_stream_conv2d_25_source_23_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_23_source_pat_fsm_5 <= _stream_conv2d_25_source_23_source_pat_fsm_5_2;
          end 
        end
        _stream_conv2d_25_source_23_source_pat_fsm_5_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_23_source_pat_fsm_5 <= _stream_conv2d_25_source_23_source_pat_fsm_5_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_24_source_pat_fsm_6_1 = 1;
  localparam _stream_conv2d_25_source_24_source_pat_fsm_6_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_24_source_pat_fsm_6 <= _stream_conv2d_25_source_24_source_pat_fsm_6_init;
    end else begin
      case(_stream_conv2d_25_source_24_source_pat_fsm_6)
        _stream_conv2d_25_source_24_source_pat_fsm_6_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_24_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_24_source_pat_fsm_6 <= _stream_conv2d_25_source_24_source_pat_fsm_6_1;
          end 
        end
        _stream_conv2d_25_source_24_source_pat_fsm_6_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_24_source_pat_fsm_6 <= _stream_conv2d_25_source_24_source_pat_fsm_6_init;
          end 
          if((_source_stream_conv2d_25_source_24_pat_count_0 == 0) && (_source_stream_conv2d_25_source_24_pat_count_1 == 0) && (_source_stream_conv2d_25_source_24_pat_count_2 == 0) && (_source_stream_conv2d_25_source_24_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_24_source_pat_fsm_6 <= _stream_conv2d_25_source_24_source_pat_fsm_6_2;
          end 
        end
        _stream_conv2d_25_source_24_source_pat_fsm_6_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_24_source_pat_fsm_6 <= _stream_conv2d_25_source_24_source_pat_fsm_6_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_25_source_pat_fsm_7_1 = 1;
  localparam _stream_conv2d_25_source_25_source_pat_fsm_7_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_25_source_pat_fsm_7 <= _stream_conv2d_25_source_25_source_pat_fsm_7_init;
    end else begin
      case(_stream_conv2d_25_source_25_source_pat_fsm_7)
        _stream_conv2d_25_source_25_source_pat_fsm_7_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_25_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_25_source_pat_fsm_7 <= _stream_conv2d_25_source_25_source_pat_fsm_7_1;
          end 
        end
        _stream_conv2d_25_source_25_source_pat_fsm_7_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_25_source_pat_fsm_7 <= _stream_conv2d_25_source_25_source_pat_fsm_7_init;
          end 
          if((_source_stream_conv2d_25_source_25_pat_count_0 == 0) && (_source_stream_conv2d_25_source_25_pat_count_1 == 0) && (_source_stream_conv2d_25_source_25_pat_count_2 == 0) && (_source_stream_conv2d_25_source_25_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_25_source_pat_fsm_7 <= _stream_conv2d_25_source_25_source_pat_fsm_7_2;
          end 
        end
        _stream_conv2d_25_source_25_source_pat_fsm_7_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_25_source_pat_fsm_7 <= _stream_conv2d_25_source_25_source_pat_fsm_7_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_26_source_pat_fsm_8_1 = 1;
  localparam _stream_conv2d_25_source_26_source_pat_fsm_8_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_26_source_pat_fsm_8 <= _stream_conv2d_25_source_26_source_pat_fsm_8_init;
    end else begin
      case(_stream_conv2d_25_source_26_source_pat_fsm_8)
        _stream_conv2d_25_source_26_source_pat_fsm_8_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_26_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_26_source_pat_fsm_8 <= _stream_conv2d_25_source_26_source_pat_fsm_8_1;
          end 
        end
        _stream_conv2d_25_source_26_source_pat_fsm_8_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_26_source_pat_fsm_8 <= _stream_conv2d_25_source_26_source_pat_fsm_8_init;
          end 
          if((_source_stream_conv2d_25_source_26_pat_count_0 == 0) && (_source_stream_conv2d_25_source_26_pat_count_1 == 0) && (_source_stream_conv2d_25_source_26_pat_count_2 == 0) && (_source_stream_conv2d_25_source_26_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_26_source_pat_fsm_8 <= _stream_conv2d_25_source_26_source_pat_fsm_8_2;
          end 
        end
        _stream_conv2d_25_source_26_source_pat_fsm_8_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_26_source_pat_fsm_8 <= _stream_conv2d_25_source_26_source_pat_fsm_8_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_27_source_pat_fsm_9_1 = 1;
  localparam _stream_conv2d_25_source_27_source_pat_fsm_9_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_27_source_pat_fsm_9 <= _stream_conv2d_25_source_27_source_pat_fsm_9_init;
    end else begin
      case(_stream_conv2d_25_source_27_source_pat_fsm_9)
        _stream_conv2d_25_source_27_source_pat_fsm_9_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_27_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_27_source_pat_fsm_9 <= _stream_conv2d_25_source_27_source_pat_fsm_9_1;
          end 
        end
        _stream_conv2d_25_source_27_source_pat_fsm_9_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_27_source_pat_fsm_9 <= _stream_conv2d_25_source_27_source_pat_fsm_9_init;
          end 
          if((_source_stream_conv2d_25_source_27_pat_count_0 == 0) && (_source_stream_conv2d_25_source_27_pat_count_1 == 0) && (_source_stream_conv2d_25_source_27_pat_count_2 == 0) && (_source_stream_conv2d_25_source_27_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_27_source_pat_fsm_9 <= _stream_conv2d_25_source_27_source_pat_fsm_9_2;
          end 
        end
        _stream_conv2d_25_source_27_source_pat_fsm_9_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_27_source_pat_fsm_9 <= _stream_conv2d_25_source_27_source_pat_fsm_9_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_28_source_pat_fsm_10_1 = 1;
  localparam _stream_conv2d_25_source_28_source_pat_fsm_10_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_28_source_pat_fsm_10 <= _stream_conv2d_25_source_28_source_pat_fsm_10_init;
    end else begin
      case(_stream_conv2d_25_source_28_source_pat_fsm_10)
        _stream_conv2d_25_source_28_source_pat_fsm_10_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_28_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_28_source_pat_fsm_10 <= _stream_conv2d_25_source_28_source_pat_fsm_10_1;
          end 
        end
        _stream_conv2d_25_source_28_source_pat_fsm_10_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_28_source_pat_fsm_10 <= _stream_conv2d_25_source_28_source_pat_fsm_10_init;
          end 
          if((_source_stream_conv2d_25_source_28_pat_count_0 == 0) && (_source_stream_conv2d_25_source_28_pat_count_1 == 0) && (_source_stream_conv2d_25_source_28_pat_count_2 == 0) && (_source_stream_conv2d_25_source_28_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_28_source_pat_fsm_10 <= _stream_conv2d_25_source_28_source_pat_fsm_10_2;
          end 
        end
        _stream_conv2d_25_source_28_source_pat_fsm_10_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_28_source_pat_fsm_10 <= _stream_conv2d_25_source_28_source_pat_fsm_10_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_29_source_pat_fsm_11_1 = 1;
  localparam _stream_conv2d_25_source_29_source_pat_fsm_11_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_29_source_pat_fsm_11 <= _stream_conv2d_25_source_29_source_pat_fsm_11_init;
    end else begin
      case(_stream_conv2d_25_source_29_source_pat_fsm_11)
        _stream_conv2d_25_source_29_source_pat_fsm_11_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_29_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_29_source_pat_fsm_11 <= _stream_conv2d_25_source_29_source_pat_fsm_11_1;
          end 
        end
        _stream_conv2d_25_source_29_source_pat_fsm_11_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_29_source_pat_fsm_11 <= _stream_conv2d_25_source_29_source_pat_fsm_11_init;
          end 
          if((_source_stream_conv2d_25_source_29_pat_count_0 == 0) && (_source_stream_conv2d_25_source_29_pat_count_1 == 0) && (_source_stream_conv2d_25_source_29_pat_count_2 == 0) && (_source_stream_conv2d_25_source_29_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_29_source_pat_fsm_11 <= _stream_conv2d_25_source_29_source_pat_fsm_11_2;
          end 
        end
        _stream_conv2d_25_source_29_source_pat_fsm_11_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_29_source_pat_fsm_11 <= _stream_conv2d_25_source_29_source_pat_fsm_11_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_30_source_pat_fsm_12_1 = 1;
  localparam _stream_conv2d_25_source_30_source_pat_fsm_12_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_30_source_pat_fsm_12 <= _stream_conv2d_25_source_30_source_pat_fsm_12_init;
    end else begin
      case(_stream_conv2d_25_source_30_source_pat_fsm_12)
        _stream_conv2d_25_source_30_source_pat_fsm_12_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_30_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_30_source_pat_fsm_12 <= _stream_conv2d_25_source_30_source_pat_fsm_12_1;
          end 
        end
        _stream_conv2d_25_source_30_source_pat_fsm_12_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_30_source_pat_fsm_12 <= _stream_conv2d_25_source_30_source_pat_fsm_12_init;
          end 
          if((_source_stream_conv2d_25_source_30_pat_count_0 == 0) && (_source_stream_conv2d_25_source_30_pat_count_1 == 0) && (_source_stream_conv2d_25_source_30_pat_count_2 == 0) && (_source_stream_conv2d_25_source_30_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_30_source_pat_fsm_12 <= _stream_conv2d_25_source_30_source_pat_fsm_12_2;
          end 
        end
        _stream_conv2d_25_source_30_source_pat_fsm_12_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_30_source_pat_fsm_12 <= _stream_conv2d_25_source_30_source_pat_fsm_12_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_31_source_pat_fsm_13_1 = 1;
  localparam _stream_conv2d_25_source_31_source_pat_fsm_13_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_31_source_pat_fsm_13 <= _stream_conv2d_25_source_31_source_pat_fsm_13_init;
    end else begin
      case(_stream_conv2d_25_source_31_source_pat_fsm_13)
        _stream_conv2d_25_source_31_source_pat_fsm_13_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_31_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_31_source_pat_fsm_13 <= _stream_conv2d_25_source_31_source_pat_fsm_13_1;
          end 
        end
        _stream_conv2d_25_source_31_source_pat_fsm_13_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_31_source_pat_fsm_13 <= _stream_conv2d_25_source_31_source_pat_fsm_13_init;
          end 
          if((_source_stream_conv2d_25_source_31_pat_count_0 == 0) && (_source_stream_conv2d_25_source_31_pat_count_1 == 0) && (_source_stream_conv2d_25_source_31_pat_count_2 == 0) && (_source_stream_conv2d_25_source_31_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_31_source_pat_fsm_13 <= _stream_conv2d_25_source_31_source_pat_fsm_13_2;
          end 
        end
        _stream_conv2d_25_source_31_source_pat_fsm_13_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_31_source_pat_fsm_13 <= _stream_conv2d_25_source_31_source_pat_fsm_13_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_32_source_pat_fsm_14_1 = 1;
  localparam _stream_conv2d_25_source_32_source_pat_fsm_14_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_32_source_pat_fsm_14 <= _stream_conv2d_25_source_32_source_pat_fsm_14_init;
    end else begin
      case(_stream_conv2d_25_source_32_source_pat_fsm_14)
        _stream_conv2d_25_source_32_source_pat_fsm_14_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_32_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_32_source_pat_fsm_14 <= _stream_conv2d_25_source_32_source_pat_fsm_14_1;
          end 
        end
        _stream_conv2d_25_source_32_source_pat_fsm_14_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_32_source_pat_fsm_14 <= _stream_conv2d_25_source_32_source_pat_fsm_14_init;
          end 
          if((_source_stream_conv2d_25_source_32_pat_count_0 == 0) && (_source_stream_conv2d_25_source_32_pat_count_1 == 0) && (_source_stream_conv2d_25_source_32_pat_count_2 == 0) && (_source_stream_conv2d_25_source_32_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_32_source_pat_fsm_14 <= _stream_conv2d_25_source_32_source_pat_fsm_14_2;
          end 
        end
        _stream_conv2d_25_source_32_source_pat_fsm_14_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_32_source_pat_fsm_14 <= _stream_conv2d_25_source_32_source_pat_fsm_14_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_33_source_pat_fsm_15_1 = 1;
  localparam _stream_conv2d_25_source_33_source_pat_fsm_15_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_33_source_pat_fsm_15 <= _stream_conv2d_25_source_33_source_pat_fsm_15_init;
    end else begin
      case(_stream_conv2d_25_source_33_source_pat_fsm_15)
        _stream_conv2d_25_source_33_source_pat_fsm_15_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_33_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_33_source_pat_fsm_15 <= _stream_conv2d_25_source_33_source_pat_fsm_15_1;
          end 
        end
        _stream_conv2d_25_source_33_source_pat_fsm_15_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_33_source_pat_fsm_15 <= _stream_conv2d_25_source_33_source_pat_fsm_15_init;
          end 
          if((_source_stream_conv2d_25_source_33_pat_count_0 == 0) && (_source_stream_conv2d_25_source_33_pat_count_1 == 0) && (_source_stream_conv2d_25_source_33_pat_count_2 == 0) && (_source_stream_conv2d_25_source_33_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_33_source_pat_fsm_15 <= _stream_conv2d_25_source_33_source_pat_fsm_15_2;
          end 
        end
        _stream_conv2d_25_source_33_source_pat_fsm_15_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_33_source_pat_fsm_15 <= _stream_conv2d_25_source_33_source_pat_fsm_15_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_34_source_pat_fsm_16_1 = 1;
  localparam _stream_conv2d_25_source_34_source_pat_fsm_16_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_34_source_pat_fsm_16 <= _stream_conv2d_25_source_34_source_pat_fsm_16_init;
    end else begin
      case(_stream_conv2d_25_source_34_source_pat_fsm_16)
        _stream_conv2d_25_source_34_source_pat_fsm_16_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_34_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_34_source_pat_fsm_16 <= _stream_conv2d_25_source_34_source_pat_fsm_16_1;
          end 
        end
        _stream_conv2d_25_source_34_source_pat_fsm_16_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_34_source_pat_fsm_16 <= _stream_conv2d_25_source_34_source_pat_fsm_16_init;
          end 
          if((_source_stream_conv2d_25_source_34_pat_count_0 == 0) && (_source_stream_conv2d_25_source_34_pat_count_1 == 0) && (_source_stream_conv2d_25_source_34_pat_count_2 == 0) && (_source_stream_conv2d_25_source_34_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_34_source_pat_fsm_16 <= _stream_conv2d_25_source_34_source_pat_fsm_16_2;
          end 
        end
        _stream_conv2d_25_source_34_source_pat_fsm_16_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_34_source_pat_fsm_16 <= _stream_conv2d_25_source_34_source_pat_fsm_16_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_35_source_pat_fsm_17_1 = 1;
  localparam _stream_conv2d_25_source_35_source_pat_fsm_17_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_35_source_pat_fsm_17 <= _stream_conv2d_25_source_35_source_pat_fsm_17_init;
    end else begin
      case(_stream_conv2d_25_source_35_source_pat_fsm_17)
        _stream_conv2d_25_source_35_source_pat_fsm_17_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_35_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_35_source_pat_fsm_17 <= _stream_conv2d_25_source_35_source_pat_fsm_17_1;
          end 
        end
        _stream_conv2d_25_source_35_source_pat_fsm_17_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_35_source_pat_fsm_17 <= _stream_conv2d_25_source_35_source_pat_fsm_17_init;
          end 
          if((_source_stream_conv2d_25_source_35_pat_count_0 == 0) && (_source_stream_conv2d_25_source_35_pat_count_1 == 0) && (_source_stream_conv2d_25_source_35_pat_count_2 == 0) && (_source_stream_conv2d_25_source_35_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_35_source_pat_fsm_17 <= _stream_conv2d_25_source_35_source_pat_fsm_17_2;
          end 
        end
        _stream_conv2d_25_source_35_source_pat_fsm_17_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_35_source_pat_fsm_17 <= _stream_conv2d_25_source_35_source_pat_fsm_17_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_36_source_pat_fsm_18_1 = 1;
  localparam _stream_conv2d_25_source_36_source_pat_fsm_18_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_36_source_pat_fsm_18 <= _stream_conv2d_25_source_36_source_pat_fsm_18_init;
    end else begin
      case(_stream_conv2d_25_source_36_source_pat_fsm_18)
        _stream_conv2d_25_source_36_source_pat_fsm_18_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_36_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_36_source_pat_fsm_18 <= _stream_conv2d_25_source_36_source_pat_fsm_18_1;
          end 
        end
        _stream_conv2d_25_source_36_source_pat_fsm_18_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_36_source_pat_fsm_18 <= _stream_conv2d_25_source_36_source_pat_fsm_18_init;
          end 
          if((_source_stream_conv2d_25_source_36_pat_count_0 == 0) && (_source_stream_conv2d_25_source_36_pat_count_1 == 0) && (_source_stream_conv2d_25_source_36_pat_count_2 == 0) && (_source_stream_conv2d_25_source_36_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_36_source_pat_fsm_18 <= _stream_conv2d_25_source_36_source_pat_fsm_18_2;
          end 
        end
        _stream_conv2d_25_source_36_source_pat_fsm_18_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_36_source_pat_fsm_18 <= _stream_conv2d_25_source_36_source_pat_fsm_18_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_source_37_source_pat_fsm_19_1 = 1;
  localparam _stream_conv2d_25_source_37_source_pat_fsm_19_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_source_37_source_pat_fsm_19 <= _stream_conv2d_25_source_37_source_pat_fsm_19_init;
    end else begin
      case(_stream_conv2d_25_source_37_source_pat_fsm_19)
        _stream_conv2d_25_source_37_source_pat_fsm_19_init: begin
          if(_stream_conv2d_25_source_start && _stream_conv2d_25_source_37_source_mode & 5'b10 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_37_source_pat_fsm_19 <= _stream_conv2d_25_source_37_source_pat_fsm_19_1;
          end 
        end
        _stream_conv2d_25_source_37_source_pat_fsm_19_1: begin
          if(_stream_conv2d_25_source_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_37_source_pat_fsm_19 <= _stream_conv2d_25_source_37_source_pat_fsm_19_init;
          end 
          if((_source_stream_conv2d_25_source_37_pat_count_0 == 0) && (_source_stream_conv2d_25_source_37_pat_count_1 == 0) && (_source_stream_conv2d_25_source_37_pat_count_2 == 0) && (_source_stream_conv2d_25_source_37_pat_count_3 == 0) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_37_source_pat_fsm_19 <= _stream_conv2d_25_source_37_source_pat_fsm_19_2;
          end 
        end
        _stream_conv2d_25_source_37_source_pat_fsm_19_2: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_source_37_source_pat_fsm_19 <= _stream_conv2d_25_source_37_source_pat_fsm_19_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_25_sink_50_sink_fsm_20_1 = 1;
  localparam _stream_conv2d_25_sink_50_sink_fsm_20_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_25_sink_50_sink_fsm_20 <= _stream_conv2d_25_sink_50_sink_fsm_20_init;
    end else begin
      case(_stream_conv2d_25_sink_50_sink_fsm_20)
        _stream_conv2d_25_sink_50_sink_fsm_20_init: begin
          if(_stream_conv2d_25_sink_start && _stream_conv2d_25_sink_50_sink_mode & 5'b1 && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_sink_50_sink_fsm_20 <= _stream_conv2d_25_sink_50_sink_fsm_20_1;
          end 
        end
        _stream_conv2d_25_sink_50_sink_fsm_20_1: begin
          if(_stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_sink_50_sink_fsm_20 <= _stream_conv2d_25_sink_50_sink_fsm_20_2;
          end 
        end
        _stream_conv2d_25_sink_50_sink_fsm_20_2: begin
          if(stream_conv2d_25_sink_51_data && (_stream_conv2d_25_sink_50_sink_count == 1) && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_sink_50_sink_fsm_20 <= _stream_conv2d_25_sink_50_sink_fsm_20_init;
          end 
          if(_stream_conv2d_25_sink_stop && _stream_conv2d_25_stream_oready) begin
            _stream_conv2d_25_sink_50_sink_fsm_20 <= _stream_conv2d_25_sink_50_sink_fsm_20_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_write_req_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_write_req_fsm <= _maxi_write_req_fsm_init;
      _maxi_write_cont <= 0;
    end else begin
      case(_maxi_write_req_fsm)
        _maxi_write_req_fsm_init: begin
          if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full) begin
            _maxi_write_req_fsm <= _maxi_write_req_fsm_1;
          end 
        end
        _maxi_write_req_fsm_1: begin
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6)) begin
            _maxi_write_cont <= 1;
          end 
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6) && (_maxi_write_global_size == 0)) begin
            _maxi_write_cont <= 0;
          end 
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6)) begin
            _maxi_write_req_fsm <= _maxi_write_req_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_write_data_fsm_1 = 1;
  localparam _maxi_write_data_fsm_2 = 2;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
    end else begin
      case(_maxi_write_data_fsm)
        _maxi_write_data_fsm_init: begin
          if(!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1)) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_1;
          end 
          if(!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2)) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_1;
          end 
          if(!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 3)) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_1;
          end 
        end
        _maxi_write_data_fsm_1: begin
          _maxi_write_data_fsm <= _maxi_write_data_fsm_2;
          _maxi_write_data_fsm <= _maxi_write_data_fsm_2;
          _maxi_write_data_fsm <= _maxi_write_data_fsm_2;
        end
        _maxi_write_data_fsm_2: begin
          if((_maxi_write_op_sel_buf == 1) && read_burst_rvalid_953 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && read_burst_rlast_954) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
          end 
          if((_maxi_write_op_sel_buf == 2) && read_burst_rvalid_1059 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && read_burst_rlast_1060) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
          end 
          if((_maxi_write_op_sel_buf == 3) && read_burst_rvalid_1199 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && read_burst_rlast_1200) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_fsm_24_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_fsm_24 <= read_burst_fsm_24_init;
      read_burst_addr_950 <= 0;
      read_burst_stride_951 <= 0;
      read_burst_length_952 <= 0;
      read_burst_rvalid_953 <= 0;
      read_burst_rlast_954 <= 0;
    end else begin
      case(read_burst_fsm_24)
        read_burst_fsm_24_init: begin
          read_burst_addr_950 <= _maxi_write_local_addr_buf;
          read_burst_stride_951 <= _maxi_write_local_stride_buf;
          read_burst_length_952 <= _maxi_write_size_buf;
          read_burst_rvalid_953 <= 0;
          read_burst_rlast_954 <= 0;
          if((_maxi_write_data_fsm == 1) && (_maxi_write_op_sel_buf == 1) && (_maxi_write_size_buf > 0)) begin
            read_burst_fsm_24 <= read_burst_fsm_24_1;
          end 
        end
        read_burst_fsm_24_1: begin
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_length_952 > 0)) begin
            read_burst_addr_950 <= read_burst_addr_950 + read_burst_stride_951;
            read_burst_length_952 <= read_burst_length_952 - 1;
            read_burst_rvalid_953 <= 1;
          end 
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_length_952 <= 1)) begin
            read_burst_rlast_954 <= 1;
          end 
          if(read_burst_rlast_954 && read_burst_rvalid_953 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_rvalid_953 <= 0;
            read_burst_rlast_954 <= 0;
          end 
          if(0) begin
            read_burst_rvalid_953 <= 0;
            read_burst_rlast_954 <= 0;
          end 
          if(read_burst_rlast_954 && read_burst_rvalid_953 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_fsm_24 <= read_burst_fsm_24_init;
          end 
          if(0) begin
            read_burst_fsm_24 <= read_burst_fsm_24_init;
          end 
        end
      endcase
    end
  end

  localparam control_max_pool_serial_27_1 = 1;
  localparam control_max_pool_serial_27_2 = 2;
  localparam control_max_pool_serial_27_3 = 3;
  localparam control_max_pool_serial_27_4 = 4;
  localparam control_max_pool_serial_27_5 = 5;
  localparam control_max_pool_serial_27_6 = 6;
  localparam control_max_pool_serial_27_7 = 7;
  localparam control_max_pool_serial_27_8 = 8;
  localparam control_max_pool_serial_27_9 = 9;
  localparam control_max_pool_serial_27_10 = 10;
  localparam control_max_pool_serial_27_11 = 11;
  localparam control_max_pool_serial_27_12 = 12;
  localparam control_max_pool_serial_27_13 = 13;
  localparam control_max_pool_serial_27_14 = 14;
  localparam control_max_pool_serial_27_15 = 15;
  localparam control_max_pool_serial_27_16 = 16;
  localparam control_max_pool_serial_27_17 = 17;
  localparam control_max_pool_serial_27_18 = 18;
  localparam control_max_pool_serial_27_19 = 19;

  always @(posedge CLK) begin
    if(RST) begin
      control_max_pool_serial_27 <= control_max_pool_serial_27_init;
      _control_max_pool_serial_27_called <= 0;
      max_pool_serial_27_act_base_offset_row <= 0;
      max_pool_serial_27_act_base_offset_bat <= 0;
      max_pool_serial_27_act_page <= 0;
      max_pool_serial_27_act_page_comp_offset <= 0;
      max_pool_serial_27_act_page_dma_offset <= 0;
      max_pool_serial_27_out_base_offset_row <= 0;
      max_pool_serial_27_out_base_offset_bat <= 0;
      max_pool_serial_27_out_page <= 0;
      max_pool_serial_27_out_page_comp_offset <= 0;
      max_pool_serial_27_out_page_dma_offset <= 0;
      max_pool_serial_27_row_count <= 0;
      max_pool_serial_27_bat_count <= 0;
      max_pool_serial_27_prev_row_count <= 0;
      max_pool_serial_27_prev_bat_count <= 0;
      max_pool_serial_27_skip_read_act <= 0;
      max_pool_serial_27_skip_comp <= 0;
      max_pool_serial_27_skip_write_out <= 0;
      max_pool_serial_27_out_count <= 0;
    end else begin
      case(control_max_pool_serial_27)
        control_max_pool_serial_27_init: begin
          if(main_fsm == 18) begin
            _control_max_pool_serial_27_called <= 1;
          end 
          if(main_fsm == 35) begin
            _control_max_pool_serial_27_called <= 1;
          end 
          if(main_fsm == 52) begin
            _control_max_pool_serial_27_called <= 1;
          end 
          if(main_fsm == 69) begin
            _control_max_pool_serial_27_called <= 1;
          end 
          if(main_fsm == 86) begin
            _control_max_pool_serial_27_called <= 1;
          end 
          if(main_fsm == 18) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_1;
          end 
          if(main_fsm == 35) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_1;
          end 
          if(main_fsm == 52) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_1;
          end 
          if(main_fsm == 69) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_1;
          end 
          if(main_fsm == 86) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_1;
          end 
        end
        control_max_pool_serial_27_1: begin
          control_max_pool_serial_27 <= control_max_pool_serial_27_2;
        end
        control_max_pool_serial_27_2: begin
          max_pool_serial_27_act_base_offset_row <= 0;
          max_pool_serial_27_act_base_offset_bat <= 0;
          max_pool_serial_27_act_page <= 0;
          max_pool_serial_27_act_page_comp_offset <= 0;
          max_pool_serial_27_act_page_dma_offset <= 0;
          max_pool_serial_27_out_base_offset_row <= 0;
          max_pool_serial_27_out_base_offset_bat <= 0;
          max_pool_serial_27_out_page <= 0;
          max_pool_serial_27_out_page_comp_offset <= 0;
          max_pool_serial_27_out_page_dma_offset <= 0;
          max_pool_serial_27_row_count <= 0;
          max_pool_serial_27_bat_count <= 0;
          max_pool_serial_27_prev_row_count <= 0;
          max_pool_serial_27_prev_bat_count <= 0;
          max_pool_serial_27_skip_read_act <= 0;
          max_pool_serial_27_skip_comp <= 0;
          max_pool_serial_27_skip_write_out <= 1;
          max_pool_serial_27_out_count <= 0;
          control_max_pool_serial_27 <= control_max_pool_serial_27_3;
        end
        control_max_pool_serial_27_3: begin
          control_max_pool_serial_27 <= control_max_pool_serial_27_4;
          if(max_pool_serial_27_skip_read_act) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_11;
          end 
        end
        control_max_pool_serial_27_4: begin
          control_max_pool_serial_27 <= control_max_pool_serial_27_5;
          if(max_pool_serial_27_dma_pad_mask_0) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_7;
          end 
        end
        control_max_pool_serial_27_5: begin
          if(_maxi_read_req_idle) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_6;
          end 
        end
        control_max_pool_serial_27_6: begin
          if(_maxi_read_idle) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_7;
          end 
        end
        control_max_pool_serial_27_7: begin
          control_max_pool_serial_27 <= control_max_pool_serial_27_8;
          if(max_pool_serial_27_dma_pad_mask_1) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_10;
          end 
        end
        control_max_pool_serial_27_8: begin
          if(_maxi_read_req_idle) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_9;
          end 
        end
        control_max_pool_serial_27_9: begin
          if(_maxi_read_idle) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_10;
          end 
        end
        control_max_pool_serial_27_10: begin
          control_max_pool_serial_27 <= control_max_pool_serial_27_11;
        end
        control_max_pool_serial_27_11: begin
          if(_maxi_write_idle) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_12;
          end 
        end
        control_max_pool_serial_27_12: begin
          if(max_pool_serial_27_comp_fsm == 0) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_13;
          end 
        end
        control_max_pool_serial_27_13: begin
          control_max_pool_serial_27 <= control_max_pool_serial_27_14;
          if(max_pool_serial_27_skip_write_out) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_17;
          end 
        end
        control_max_pool_serial_27_14: begin
          if(max_pool_serial_27_comp_count >= max_pool_serial_27_out_count + cparam_max_pool_serial_27_out_write_size) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_15;
          end 
        end
        control_max_pool_serial_27_15: begin
          if(_maxi_write_req_idle) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_16;
          end 
        end
        control_max_pool_serial_27_16: begin
          max_pool_serial_27_out_count <= max_pool_serial_27_out_count + cparam_max_pool_serial_27_out_write_size;
          control_max_pool_serial_27 <= control_max_pool_serial_27_17;
        end
        control_max_pool_serial_27_17: begin
          max_pool_serial_27_act_base_offset_row <= max_pool_serial_27_act_base_offset_row + cparam_max_pool_serial_27_act_row_step;
          if(max_pool_serial_27_row_count >= cparam_max_pool_serial_27_max_row_count) begin
            max_pool_serial_27_act_base_offset_row <= 0;
            max_pool_serial_27_act_base_offset_bat <= max_pool_serial_27_act_base_offset_bat + cparam_max_pool_serial_27_act_bat_step;
          end 
          if((max_pool_serial_27_row_count >= cparam_max_pool_serial_27_max_row_count) && (max_pool_serial_27_bat_count >= cparam_max_pool_serial_27_max_bat_count)) begin
            max_pool_serial_27_act_base_offset_bat <= 0;
          end 
          max_pool_serial_27_row_count <= max_pool_serial_27_row_count + cparam_max_pool_serial_27_stride_row;
          if(max_pool_serial_27_row_count >= cparam_max_pool_serial_27_max_row_count) begin
            max_pool_serial_27_row_count <= 0;
            max_pool_serial_27_bat_count <= max_pool_serial_27_bat_count + 1;
          end 
          if((max_pool_serial_27_row_count >= cparam_max_pool_serial_27_max_row_count) && (max_pool_serial_27_bat_count >= cparam_max_pool_serial_27_max_bat_count)) begin
            max_pool_serial_27_bat_count <= 0;
          end 
          if(!max_pool_serial_27_act_page) begin
            max_pool_serial_27_act_page_comp_offset <= 16384;
            max_pool_serial_27_act_page_dma_offset <= 16384;
            max_pool_serial_27_act_page <= 1;
          end 
          if(max_pool_serial_27_act_page) begin
            max_pool_serial_27_act_page_comp_offset <= 0;
            max_pool_serial_27_act_page_dma_offset <= 0;
            max_pool_serial_27_act_page <= 0;
          end 
          if(!max_pool_serial_27_skip_write_out) begin
            max_pool_serial_27_out_base_offset_row <= max_pool_serial_27_out_base_offset_row + cparam_max_pool_serial_27_out_row_step;
          end 
          if(!max_pool_serial_27_skip_write_out && (max_pool_serial_27_prev_row_count >= cparam_max_pool_serial_27_max_row_count)) begin
            max_pool_serial_27_out_base_offset_row <= 0;
            max_pool_serial_27_out_base_offset_bat <= max_pool_serial_27_out_base_offset_bat + cparam_max_pool_serial_27_out_bat_step;
          end 
          if(!max_pool_serial_27_skip_write_out && (max_pool_serial_27_prev_row_count >= cparam_max_pool_serial_27_max_row_count) && (max_pool_serial_27_prev_bat_count >= cparam_max_pool_serial_27_max_bat_count)) begin
            max_pool_serial_27_out_base_offset_bat <= 0;
          end 
          if(!max_pool_serial_27_out_page) begin
            max_pool_serial_27_out_page_comp_offset <= 4096;
            max_pool_serial_27_out_page_dma_offset <= 0;
            max_pool_serial_27_out_page <= 1;
          end 
          if(max_pool_serial_27_out_page) begin
            max_pool_serial_27_out_page_comp_offset <= 0;
            max_pool_serial_27_out_page_dma_offset <= 4096;
            max_pool_serial_27_out_page <= 0;
          end 
          max_pool_serial_27_prev_row_count <= max_pool_serial_27_row_count;
          max_pool_serial_27_prev_bat_count <= max_pool_serial_27_bat_count;
          if((max_pool_serial_27_row_count >= cparam_max_pool_serial_27_max_row_count) && (max_pool_serial_27_bat_count >= cparam_max_pool_serial_27_max_bat_count)) begin
            max_pool_serial_27_skip_read_act <= 1;
          end 
          if((max_pool_serial_27_row_count >= cparam_max_pool_serial_27_max_row_count) && (max_pool_serial_27_bat_count >= cparam_max_pool_serial_27_max_bat_count)) begin
            max_pool_serial_27_skip_comp <= 1;
          end 
          if(max_pool_serial_27_skip_write_out && (max_pool_serial_27_prev_row_count == 0) && (max_pool_serial_27_prev_bat_count == 0)) begin
            max_pool_serial_27_skip_write_out <= 0;
          end 
          control_max_pool_serial_27 <= control_max_pool_serial_27_3;
          if(!max_pool_serial_27_skip_write_out && (max_pool_serial_27_prev_row_count >= cparam_max_pool_serial_27_max_row_count) && (max_pool_serial_27_prev_bat_count >= cparam_max_pool_serial_27_max_bat_count)) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_18;
          end 
        end
        control_max_pool_serial_27_18: begin
          if(_maxi_write_idle && !_maxi_has_outstanding_write) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_19;
          end 
        end
        control_max_pool_serial_27_19: begin
          if(main_fsm == 21) begin
            _control_max_pool_serial_27_called <= 0;
          end 
          if(main_fsm == 38) begin
            _control_max_pool_serial_27_called <= 0;
          end 
          if(main_fsm == 55) begin
            _control_max_pool_serial_27_called <= 0;
          end 
          if(main_fsm == 72) begin
            _control_max_pool_serial_27_called <= 0;
          end 
          if(main_fsm == 89) begin
            _control_max_pool_serial_27_called <= 0;
          end 
          if(main_fsm == 21) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_init;
          end 
          if(main_fsm == 38) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_init;
          end 
          if(main_fsm == 55) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_init;
          end 
          if(main_fsm == 72) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_init;
          end 
          if(main_fsm == 89) begin
            control_max_pool_serial_27 <= control_max_pool_serial_27_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_25_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_25 <= write_burst_fsm_25_init;
      write_burst_addr_960 <= 0;
      write_burst_stride_961 <= 0;
      write_burst_length_962 <= 0;
      write_burst_done_963 <= 0;
    end else begin
      case(write_burst_fsm_25)
        write_burst_fsm_25_init: begin
          write_burst_addr_960 <= _maxi_read_local_addr_buf;
          write_burst_stride_961 <= _maxi_read_local_stride_buf;
          write_burst_length_962 <= _maxi_read_local_size_buf;
          write_burst_done_963 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 7) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_25 <= write_burst_fsm_25_1;
          end 
        end
        write_burst_fsm_25_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_addr_960 <= write_burst_addr_960 + write_burst_stride_961;
            write_burst_length_962 <= write_burst_length_962 - 1;
            write_burst_done_963 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_962 <= 1)) begin
            write_burst_done_963 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_done_963 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_962 <= 1)) begin
            write_burst_fsm_25 <= write_burst_fsm_25_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_fsm_25 <= write_burst_fsm_25_init;
          end 
          if(0) begin
            write_burst_fsm_25 <= write_burst_fsm_25_init;
          end 
        end
      endcase
    end
  end

  localparam max_pool_serial_27_comp_fsm_1 = 1;
  localparam max_pool_serial_27_comp_fsm_2 = 2;
  localparam max_pool_serial_27_comp_fsm_3 = 3;
  localparam max_pool_serial_27_comp_fsm_4 = 4;
  localparam max_pool_serial_27_comp_fsm_5 = 5;
  localparam max_pool_serial_27_comp_fsm_6 = 6;
  localparam max_pool_serial_27_comp_fsm_7 = 7;

  always @(posedge CLK) begin
    if(RST) begin
      max_pool_serial_27_comp_fsm <= max_pool_serial_27_comp_fsm_init;
      max_pool_serial_27_stream_act_local <= 0;
      max_pool_serial_27_stream_out_local <= 0;
      max_pool_serial_27_col_count <= 0;
      max_pool_serial_27_act_page_comp_offset_buf <= 0;
      max_pool_serial_27_out_page_comp_offset_buf <= 0;
      max_pool_serial_27_row_count_buf <= 0;
      max_pool_serial_27_stream_pad_masks <= 0;
      max_pool_serial_27_comp_count <= 0;
    end else begin
      if(control_max_pool_serial_27 == 2) begin
        max_pool_serial_27_comp_count <= 0;
      end 
      if(_stream_max_pool_serial_27_sink_stop) begin
        max_pool_serial_27_comp_count <= max_pool_serial_27_comp_count + cparam_max_pool_serial_27_inc_out_laddr;
      end 
      case(max_pool_serial_27_comp_fsm)
        max_pool_serial_27_comp_fsm_init: begin
          if((control_max_pool_serial_27 == 12) && !max_pool_serial_27_skip_comp) begin
            max_pool_serial_27_comp_fsm <= max_pool_serial_27_comp_fsm_1;
          end 
        end
        max_pool_serial_27_comp_fsm_1: begin
          max_pool_serial_27_stream_act_local <= cparam_max_pool_serial_27_local_pad_offset;
          max_pool_serial_27_stream_out_local <= 0;
          max_pool_serial_27_col_count <= 0;
          max_pool_serial_27_act_page_comp_offset_buf <= max_pool_serial_27_act_page_comp_offset;
          max_pool_serial_27_out_page_comp_offset_buf <= max_pool_serial_27_out_page_comp_offset;
          max_pool_serial_27_row_count_buf <= max_pool_serial_27_row_count;
          max_pool_serial_27_comp_fsm <= max_pool_serial_27_comp_fsm_2;
        end
        max_pool_serial_27_comp_fsm_2: begin
          max_pool_serial_27_stream_pad_masks <= { max_pool_serial_27_stream_pad_mask_1_1, max_pool_serial_27_stream_pad_mask_1_0, max_pool_serial_27_stream_pad_mask_0_1, max_pool_serial_27_stream_pad_mask_0_0 };
          max_pool_serial_27_comp_fsm <= max_pool_serial_27_comp_fsm_3;
        end
        max_pool_serial_27_comp_fsm_3: begin
          if(!_stream_max_pool_serial_27_source_busy) begin
            max_pool_serial_27_comp_fsm <= max_pool_serial_27_comp_fsm_4;
          end 
        end
        max_pool_serial_27_comp_fsm_4: begin
          max_pool_serial_27_comp_fsm <= max_pool_serial_27_comp_fsm_5;
          max_pool_serial_27_comp_fsm <= max_pool_serial_27_comp_fsm_5;
          max_pool_serial_27_comp_fsm <= max_pool_serial_27_comp_fsm_5;
          if(_stream_max_pool_serial_27_stream_oready) begin
            max_pool_serial_27_comp_fsm <= max_pool_serial_27_comp_fsm_5;
          end 
        end
        max_pool_serial_27_comp_fsm_5: begin
          max_pool_serial_27_comp_fsm <= max_pool_serial_27_comp_fsm_6;
        end
        max_pool_serial_27_comp_fsm_6: begin
          if(_stream_max_pool_serial_27_busy) begin
            max_pool_serial_27_comp_fsm <= max_pool_serial_27_comp_fsm_7;
          end 
        end
        max_pool_serial_27_comp_fsm_7: begin
          max_pool_serial_27_stream_act_local <= max_pool_serial_27_stream_act_local + cparam_max_pool_serial_27_inc_act_laddr;
          if(max_pool_serial_27_col_count >= cparam_max_pool_serial_27_max_col_count) begin
            max_pool_serial_27_stream_act_local <= cparam_max_pool_serial_27_local_pad_offset;
          end 
          max_pool_serial_27_stream_out_local <= max_pool_serial_27_stream_out_local + cparam_max_pool_serial_27_inc_out_laddr;
          if(max_pool_serial_27_col_count >= cparam_max_pool_serial_27_max_col_count) begin
            max_pool_serial_27_stream_out_local <= 0;
          end 
          max_pool_serial_27_col_count <= max_pool_serial_27_col_count + cparam_max_pool_serial_27_stride_col;
          if(max_pool_serial_27_col_count >= cparam_max_pool_serial_27_max_col_count) begin
            max_pool_serial_27_col_count <= 0;
          end 
          max_pool_serial_27_comp_fsm <= max_pool_serial_27_comp_fsm_2;
          if(max_pool_serial_27_col_count >= cparam_max_pool_serial_27_max_col_count) begin
            max_pool_serial_27_comp_fsm <= max_pool_serial_27_comp_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_max_pool_serial_27_source_1_source_pat_fsm_0_1 = 1;
  localparam _stream_max_pool_serial_27_source_1_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_27_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_27_source_1_source_pat_fsm_0_init;
    end else begin
      case(_stream_max_pool_serial_27_source_1_source_pat_fsm_0)
        _stream_max_pool_serial_27_source_1_source_pat_fsm_0_init: begin
          if(_stream_max_pool_serial_27_source_start && _stream_max_pool_serial_27_source_1_source_mode & 5'b10 && _stream_max_pool_serial_27_stream_oready) begin
            _stream_max_pool_serial_27_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_27_source_1_source_pat_fsm_0_1;
          end 
        end
        _stream_max_pool_serial_27_source_1_source_pat_fsm_0_1: begin
          if(_stream_max_pool_serial_27_source_stop && _stream_max_pool_serial_27_stream_oready) begin
            _stream_max_pool_serial_27_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_27_source_1_source_pat_fsm_0_init;
          end 
          if((_source_stream_max_pool_serial_27_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_27_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_27_source_1_pat_count_2 == 0) && (_source_stream_max_pool_serial_27_source_1_pat_count_3 == 0) && _stream_max_pool_serial_27_stream_oready) begin
            _stream_max_pool_serial_27_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_27_source_1_source_pat_fsm_0_2;
          end 
        end
        _stream_max_pool_serial_27_source_1_source_pat_fsm_0_2: begin
          if(_stream_max_pool_serial_27_stream_oready) begin
            _stream_max_pool_serial_27_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_27_source_1_source_pat_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_max_pool_serial_27_sink_5_sink_fsm_1_1 = 1;
  localparam _stream_max_pool_serial_27_sink_5_sink_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_27_sink_5_sink_fsm_1 <= _stream_max_pool_serial_27_sink_5_sink_fsm_1_init;
    end else begin
      case(_stream_max_pool_serial_27_sink_5_sink_fsm_1)
        _stream_max_pool_serial_27_sink_5_sink_fsm_1_init: begin
          if(_stream_max_pool_serial_27_sink_start && _stream_max_pool_serial_27_sink_5_sink_mode & 5'b1 && _stream_max_pool_serial_27_stream_oready) begin
            _stream_max_pool_serial_27_sink_5_sink_fsm_1 <= _stream_max_pool_serial_27_sink_5_sink_fsm_1_1;
          end 
        end
        _stream_max_pool_serial_27_sink_5_sink_fsm_1_1: begin
          if(_stream_max_pool_serial_27_stream_oready) begin
            _stream_max_pool_serial_27_sink_5_sink_fsm_1 <= _stream_max_pool_serial_27_sink_5_sink_fsm_1_2;
          end 
        end
        _stream_max_pool_serial_27_sink_5_sink_fsm_1_2: begin
          if(stream_max_pool_serial_27_sink_6_data && (_stream_max_pool_serial_27_sink_5_sink_count == 1) && _stream_max_pool_serial_27_stream_oready) begin
            _stream_max_pool_serial_27_sink_5_sink_fsm_1 <= _stream_max_pool_serial_27_sink_5_sink_fsm_1_init;
          end 
          if(_stream_max_pool_serial_27_sink_stop && _stream_max_pool_serial_27_stream_oready) begin
            _stream_max_pool_serial_27_sink_5_sink_fsm_1 <= _stream_max_pool_serial_27_sink_5_sink_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_fsm_26_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_fsm_26 <= read_burst_fsm_26_init;
      read_burst_addr_1056 <= 0;
      read_burst_stride_1057 <= 0;
      read_burst_length_1058 <= 0;
      read_burst_rvalid_1059 <= 0;
      read_burst_rlast_1060 <= 0;
    end else begin
      case(read_burst_fsm_26)
        read_burst_fsm_26_init: begin
          read_burst_addr_1056 <= _maxi_write_local_addr_buf;
          read_burst_stride_1057 <= _maxi_write_local_stride_buf;
          read_burst_length_1058 <= _maxi_write_size_buf;
          read_burst_rvalid_1059 <= 0;
          read_burst_rlast_1060 <= 0;
          if((_maxi_write_data_fsm == 1) && (_maxi_write_op_sel_buf == 2) && (_maxi_write_size_buf > 0)) begin
            read_burst_fsm_26 <= read_burst_fsm_26_1;
          end 
        end
        read_burst_fsm_26_1: begin
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_length_1058 > 0)) begin
            read_burst_addr_1056 <= read_burst_addr_1056 + read_burst_stride_1057;
            read_burst_length_1058 <= read_burst_length_1058 - 1;
            read_burst_rvalid_1059 <= 1;
          end 
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_length_1058 <= 1)) begin
            read_burst_rlast_1060 <= 1;
          end 
          if(read_burst_rlast_1060 && read_burst_rvalid_1059 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_rvalid_1059 <= 0;
            read_burst_rlast_1060 <= 0;
          end 
          if(0) begin
            read_burst_rvalid_1059 <= 0;
            read_burst_rlast_1060 <= 0;
          end 
          if(read_burst_rlast_1060 && read_burst_rvalid_1059 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_fsm_26 <= read_burst_fsm_26_init;
          end 
          if(0) begin
            read_burst_fsm_26 <= read_burst_fsm_26_init;
          end 
        end
      endcase
    end
  end

  localparam control_max_pool_47_1 = 1;
  localparam control_max_pool_47_2 = 2;
  localparam control_max_pool_47_3 = 3;
  localparam control_max_pool_47_4 = 4;
  localparam control_max_pool_47_5 = 5;
  localparam control_max_pool_47_6 = 6;
  localparam control_max_pool_47_7 = 7;
  localparam control_max_pool_47_8 = 8;
  localparam control_max_pool_47_9 = 9;
  localparam control_max_pool_47_10 = 10;
  localparam control_max_pool_47_11 = 11;
  localparam control_max_pool_47_12 = 12;
  localparam control_max_pool_47_13 = 13;
  localparam control_max_pool_47_14 = 14;
  localparam control_max_pool_47_15 = 15;
  localparam control_max_pool_47_16 = 16;
  localparam control_max_pool_47_17 = 17;
  localparam control_max_pool_47_18 = 18;
  localparam control_max_pool_47_19 = 19;

  always @(posedge CLK) begin
    if(RST) begin
      control_max_pool_47 <= control_max_pool_47_init;
      _control_max_pool_47_called <= 0;
      max_pool_47_act_base_offset_row <= 0;
      max_pool_47_act_base_offset_bat <= 0;
      max_pool_47_dma_flag_0 <= 0;
      max_pool_47_dma_flag_1 <= 0;
      max_pool_47_act_page_0 <= 0;
      max_pool_47_act_page_1 <= 0;
      max_pool_47_act_page_comp_offset_0 <= 0;
      max_pool_47_act_page_comp_offset_1 <= 0;
      max_pool_47_act_page_dma_offset_0 <= 0;
      max_pool_47_act_page_dma_offset_1 <= 0;
      max_pool_47_out_base_offset_row <= 0;
      max_pool_47_out_base_offset_bat <= 0;
      max_pool_47_out_page <= 0;
      max_pool_47_out_page_comp_offset <= 0;
      max_pool_47_out_page_dma_offset <= 0;
      max_pool_47_row_count <= 0;
      max_pool_47_bat_count <= 0;
      max_pool_47_row_select <= 0;
      max_pool_47_prev_row_count <= 0;
      max_pool_47_prev_bat_count <= 0;
      max_pool_47_prev_row_select <= 0;
      max_pool_47_skip_read_act <= 0;
      max_pool_47_skip_comp <= 0;
      max_pool_47_skip_write_out <= 0;
      max_pool_47_out_count <= 0;
    end else begin
      case(control_max_pool_47)
        control_max_pool_47_init: begin
          if(main_fsm == 102) begin
            _control_max_pool_47_called <= 1;
          end 
          if(main_fsm == 102) begin
            control_max_pool_47 <= control_max_pool_47_1;
          end 
        end
        control_max_pool_47_1: begin
          control_max_pool_47 <= control_max_pool_47_2;
        end
        control_max_pool_47_2: begin
          max_pool_47_act_base_offset_row <= 0;
          max_pool_47_act_base_offset_bat <= 0;
          max_pool_47_dma_flag_0 <= 1;
          max_pool_47_dma_flag_1 <= 1;
          max_pool_47_act_page_0 <= 0;
          max_pool_47_act_page_1 <= 0;
          max_pool_47_act_page_comp_offset_0 <= 0;
          max_pool_47_act_page_comp_offset_1 <= 0;
          max_pool_47_act_page_dma_offset_0 <= 0;
          max_pool_47_act_page_dma_offset_1 <= 0;
          max_pool_47_out_base_offset_row <= 0;
          max_pool_47_out_base_offset_bat <= 0;
          max_pool_47_out_page <= 0;
          max_pool_47_out_page_comp_offset <= 0;
          max_pool_47_out_page_dma_offset <= 0;
          max_pool_47_row_count <= 0;
          max_pool_47_bat_count <= 0;
          max_pool_47_row_select <= 0;
          max_pool_47_prev_row_count <= 0;
          max_pool_47_prev_bat_count <= 0;
          max_pool_47_prev_row_select <= 0;
          max_pool_47_skip_read_act <= 0;
          max_pool_47_skip_comp <= 0;
          max_pool_47_skip_write_out <= 1;
          max_pool_47_out_count <= 0;
          control_max_pool_47 <= control_max_pool_47_3;
        end
        control_max_pool_47_3: begin
          control_max_pool_47 <= control_max_pool_47_4;
          if(max_pool_47_skip_read_act) begin
            control_max_pool_47 <= control_max_pool_47_11;
          end 
        end
        control_max_pool_47_4: begin
          control_max_pool_47 <= control_max_pool_47_5;
          if(max_pool_47_mux_dma_pad_mask_0 || !max_pool_47_mux_dma_flag_0) begin
            control_max_pool_47 <= control_max_pool_47_7;
          end 
        end
        control_max_pool_47_5: begin
          if(_maxi_read_req_idle) begin
            control_max_pool_47 <= control_max_pool_47_6;
          end 
        end
        control_max_pool_47_6: begin
          if(_maxi_read_idle) begin
            control_max_pool_47 <= control_max_pool_47_7;
          end 
        end
        control_max_pool_47_7: begin
          control_max_pool_47 <= control_max_pool_47_8;
          if(max_pool_47_mux_dma_pad_mask_1 || !max_pool_47_mux_dma_flag_1) begin
            control_max_pool_47 <= control_max_pool_47_10;
          end 
        end
        control_max_pool_47_8: begin
          if(_maxi_read_req_idle) begin
            control_max_pool_47 <= control_max_pool_47_9;
          end 
        end
        control_max_pool_47_9: begin
          if(_maxi_read_idle) begin
            control_max_pool_47 <= control_max_pool_47_10;
          end 
        end
        control_max_pool_47_10: begin
          control_max_pool_47 <= control_max_pool_47_11;
        end
        control_max_pool_47_11: begin
          if(_maxi_write_idle) begin
            control_max_pool_47 <= control_max_pool_47_12;
          end 
        end
        control_max_pool_47_12: begin
          if(max_pool_47_comp_fsm == 0) begin
            control_max_pool_47 <= control_max_pool_47_13;
          end 
        end
        control_max_pool_47_13: begin
          control_max_pool_47 <= control_max_pool_47_14;
          if(max_pool_47_skip_write_out) begin
            control_max_pool_47 <= control_max_pool_47_17;
          end 
        end
        control_max_pool_47_14: begin
          if(max_pool_47_comp_count >= max_pool_47_out_count + cparam_max_pool_47_out_write_size) begin
            control_max_pool_47 <= control_max_pool_47_15;
          end 
        end
        control_max_pool_47_15: begin
          if(_maxi_write_req_idle) begin
            control_max_pool_47 <= control_max_pool_47_16;
          end 
        end
        control_max_pool_47_16: begin
          max_pool_47_out_count <= max_pool_47_out_count + cparam_max_pool_47_out_write_size;
          control_max_pool_47 <= control_max_pool_47_17;
        end
        control_max_pool_47_17: begin
          max_pool_47_act_base_offset_row <= max_pool_47_act_base_offset_row + cparam_max_pool_47_act_row_step;
          if(max_pool_47_row_count >= cparam_max_pool_47_max_row_count) begin
            max_pool_47_act_base_offset_row <= 0;
            max_pool_47_act_base_offset_bat <= max_pool_47_act_base_offset_bat + cparam_max_pool_47_act_bat_step;
          end 
          if((max_pool_47_row_count >= cparam_max_pool_47_max_row_count) && (max_pool_47_bat_count >= cparam_max_pool_47_max_bat_count)) begin
            max_pool_47_act_base_offset_bat <= 0;
          end 
          max_pool_47_dma_flag_0 <= cparam_max_pool_47_dma_flag_conds_0;
          if(max_pool_47_row_count >= cparam_max_pool_47_max_row_count) begin
            max_pool_47_dma_flag_0 <= 1;
          end 
          max_pool_47_dma_flag_1 <= cparam_max_pool_47_dma_flag_conds_1;
          if(max_pool_47_row_count >= cparam_max_pool_47_max_row_count) begin
            max_pool_47_dma_flag_1 <= 1;
          end 
          max_pool_47_row_count <= max_pool_47_row_count + cparam_max_pool_47_stride_row;
          if(max_pool_47_row_count >= cparam_max_pool_47_max_row_count) begin
            max_pool_47_row_count <= 0;
            max_pool_47_bat_count <= max_pool_47_bat_count + 1;
          end 
          if((max_pool_47_row_count >= cparam_max_pool_47_max_row_count) && (max_pool_47_bat_count >= cparam_max_pool_47_max_bat_count)) begin
            max_pool_47_bat_count <= 0;
          end 
          if(cparam_max_pool_47_stride_row < 2) begin
            max_pool_47_row_select <= max_pool_47_row_select + cparam_max_pool_47_stride_row;
            max_pool_47_prev_row_select <= max_pool_47_row_select;
          end 
          if((cparam_max_pool_47_stride_row < 2) && (max_pool_47_row_select + cparam_max_pool_47_stride_row >= 2)) begin
            max_pool_47_row_select <= max_pool_47_row_select - (2 - cparam_max_pool_47_stride_row);
            max_pool_47_prev_row_select <= max_pool_47_row_select;
          end 
          if(!(cparam_max_pool_47_stride_row < 2)) begin
            max_pool_47_row_select <= 0;
            max_pool_47_prev_row_select <= 0;
          end 
          if(max_pool_47_row_count >= cparam_max_pool_47_max_row_count) begin
            max_pool_47_row_select <= 0;
            max_pool_47_prev_row_select <= 0;
          end 
          if(!max_pool_47_act_page_0 && max_pool_47_mux_next_dma_flag_0) begin
            max_pool_47_act_page_comp_offset_0 <= 4096;
            max_pool_47_act_page_dma_offset_0 <= 4096;
            max_pool_47_act_page_0 <= 1;
          end 
          if(max_pool_47_act_page_0 && max_pool_47_mux_next_dma_flag_0) begin
            max_pool_47_act_page_comp_offset_0 <= 0;
            max_pool_47_act_page_dma_offset_0 <= 0;
            max_pool_47_act_page_0 <= 0;
          end 
          if(!max_pool_47_act_page_1 && max_pool_47_mux_next_dma_flag_1) begin
            max_pool_47_act_page_comp_offset_1 <= 4096;
            max_pool_47_act_page_dma_offset_1 <= 4096;
            max_pool_47_act_page_1 <= 1;
          end 
          if(max_pool_47_act_page_1 && max_pool_47_mux_next_dma_flag_1) begin
            max_pool_47_act_page_comp_offset_1 <= 0;
            max_pool_47_act_page_dma_offset_1 <= 0;
            max_pool_47_act_page_1 <= 0;
          end 
          if(!max_pool_47_skip_write_out) begin
            max_pool_47_out_base_offset_row <= max_pool_47_out_base_offset_row + cparam_max_pool_47_out_row_step;
          end 
          if(!max_pool_47_skip_write_out && (max_pool_47_prev_row_count >= cparam_max_pool_47_max_row_count)) begin
            max_pool_47_out_base_offset_row <= 0;
            max_pool_47_out_base_offset_bat <= max_pool_47_out_base_offset_bat + cparam_max_pool_47_out_bat_step;
          end 
          if(!max_pool_47_skip_write_out && (max_pool_47_prev_row_count >= cparam_max_pool_47_max_row_count) && (max_pool_47_prev_bat_count >= cparam_max_pool_47_max_bat_count)) begin
            max_pool_47_out_base_offset_bat <= 0;
          end 
          if(!max_pool_47_out_page) begin
            max_pool_47_out_page_comp_offset <= 8192;
            max_pool_47_out_page_dma_offset <= 0;
            max_pool_47_out_page <= 1;
          end 
          if(max_pool_47_out_page) begin
            max_pool_47_out_page_comp_offset <= 0;
            max_pool_47_out_page_dma_offset <= 8192;
            max_pool_47_out_page <= 0;
          end 
          max_pool_47_prev_row_count <= max_pool_47_row_count;
          max_pool_47_prev_bat_count <= max_pool_47_bat_count;
          if((max_pool_47_row_count >= cparam_max_pool_47_max_row_count) && (max_pool_47_bat_count >= cparam_max_pool_47_max_bat_count)) begin
            max_pool_47_skip_read_act <= 1;
          end 
          if((max_pool_47_row_count >= cparam_max_pool_47_max_row_count) && (max_pool_47_bat_count >= cparam_max_pool_47_max_bat_count)) begin
            max_pool_47_skip_comp <= 1;
          end 
          if(max_pool_47_skip_write_out && (max_pool_47_prev_row_count == 0) && (max_pool_47_prev_bat_count == 0)) begin
            max_pool_47_skip_write_out <= 0;
          end 
          control_max_pool_47 <= control_max_pool_47_3;
          if(!max_pool_47_skip_write_out && (max_pool_47_prev_row_count >= cparam_max_pool_47_max_row_count) && (max_pool_47_prev_bat_count >= cparam_max_pool_47_max_bat_count)) begin
            control_max_pool_47 <= control_max_pool_47_18;
          end 
        end
        control_max_pool_47_18: begin
          if(_maxi_write_idle && !_maxi_has_outstanding_write) begin
            control_max_pool_47 <= control_max_pool_47_19;
          end 
        end
        control_max_pool_47_19: begin
          if(main_fsm == 105) begin
            _control_max_pool_47_called <= 0;
          end 
          if(main_fsm == 105) begin
            control_max_pool_47 <= control_max_pool_47_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_27_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_27 <= write_burst_fsm_27_init;
      write_burst_addr_1068 <= 0;
      write_burst_stride_1069 <= 0;
      write_burst_length_1070 <= 0;
      write_burst_done_1071 <= 0;
    end else begin
      case(write_burst_fsm_27)
        write_burst_fsm_27_init: begin
          write_burst_addr_1068 <= _maxi_read_local_addr_buf;
          write_burst_stride_1069 <= _maxi_read_local_stride_buf;
          write_burst_length_1070 <= _maxi_read_local_size_buf;
          write_burst_done_1071 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 8) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_27 <= write_burst_fsm_27_1;
          end 
        end
        write_burst_fsm_27_1: begin
          if(write_burst_block_ram_wvalid_1066) begin
            write_burst_addr_1068 <= write_burst_addr_1068 + write_burst_stride_1069;
            write_burst_length_1070 <= write_burst_length_1070 - 1;
            write_burst_done_1071 <= 0;
          end 
          if(write_burst_block_ram_wvalid_1066 && (write_burst_length_1070 <= 1)) begin
            write_burst_done_1071 <= 1;
          end 
          if(write_burst_block_ram_wvalid_1066 && 0) begin
            write_burst_done_1071 <= 1;
          end 
          if(write_burst_block_ram_wvalid_1066 && (write_burst_length_1070 <= 1)) begin
            write_burst_fsm_27 <= write_burst_fsm_27_init;
          end 
          if(write_burst_block_ram_wvalid_1066 && 0) begin
            write_burst_fsm_27 <= write_burst_fsm_27_init;
          end 
          if(write_burst_block_ram_wquit_1067) begin
            write_burst_fsm_27 <= write_burst_fsm_27_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_28_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_28 <= write_burst_fsm_28_init;
      write_burst_addr_1074 <= 0;
      write_burst_stride_1075 <= 0;
      write_burst_length_1076 <= 0;
      write_burst_done_1077 <= 0;
    end else begin
      case(write_burst_fsm_28)
        write_burst_fsm_28_init: begin
          write_burst_addr_1074 <= _maxi_read_local_addr_buf;
          write_burst_stride_1075 <= _maxi_read_local_stride_buf;
          write_burst_length_1076 <= _maxi_read_local_size_buf;
          write_burst_done_1077 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 8) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_28 <= write_burst_fsm_28_1;
          end 
        end
        write_burst_fsm_28_1: begin
          if(write_burst_block_ram_wvalid_1072) begin
            write_burst_addr_1074 <= write_burst_addr_1074 + write_burst_stride_1075;
            write_burst_length_1076 <= write_burst_length_1076 - 1;
            write_burst_done_1077 <= 0;
          end 
          if(write_burst_block_ram_wvalid_1072 && (write_burst_length_1076 <= 1)) begin
            write_burst_done_1077 <= 1;
          end 
          if(write_burst_block_ram_wvalid_1072 && 0) begin
            write_burst_done_1077 <= 1;
          end 
          if(write_burst_block_ram_wvalid_1072 && (write_burst_length_1076 <= 1)) begin
            write_burst_fsm_28 <= write_burst_fsm_28_init;
          end 
          if(write_burst_block_ram_wvalid_1072 && 0) begin
            write_burst_fsm_28 <= write_burst_fsm_28_init;
          end 
          if(write_burst_block_ram_wquit_1073) begin
            write_burst_fsm_28 <= write_burst_fsm_28_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_29_1 = 1;
  localparam write_burst_block_fsm_29_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_29 <= write_burst_block_fsm_29_init;
      write_burst_block_length_1078 <= 0;
      write_burst_block_blocksize_1079 <= 0;
      write_burst_block_done_1080 <= 0;
      write_burst_block_count_1081 <= 0;
    end else begin
      case(write_burst_block_fsm_29)
        write_burst_block_fsm_29_init: begin
          write_burst_block_length_1078 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_1079 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_1080 <= 0;
          write_burst_block_count_1081 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 8) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_29 <= write_burst_block_fsm_29_1;
          end 
        end
        write_burst_block_fsm_29_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_1078 <= write_burst_block_length_1078 - 1;
            write_burst_block_done_1080 <= 0;
            write_burst_block_count_1081 <= write_burst_block_count_1081 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_1078 <= 1)) begin
            write_burst_block_done_1080 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_1080 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_1081 == write_burst_block_blocksize_1079 - 1)) begin
            write_burst_block_count_1081 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_1081 == write_burst_block_blocksize_1079 - 1)) begin
            write_burst_block_fsm_29 <= write_burst_block_fsm_29_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_1078 <= 1)) begin
            write_burst_block_fsm_29 <= write_burst_block_fsm_29_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_29 <= write_burst_block_fsm_29_init;
          end 
          if(0) begin
            write_burst_block_fsm_29 <= write_burst_block_fsm_29_init;
          end 
        end
        write_burst_block_fsm_29_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_1078 <= write_burst_block_length_1078 - 1;
            write_burst_block_done_1080 <= 0;
            write_burst_block_count_1081 <= write_burst_block_count_1081 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_1078 <= 1)) begin
            write_burst_block_done_1080 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_1080 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_1081 == write_burst_block_blocksize_1079 - 1)) begin
            write_burst_block_count_1081 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_1081 == write_burst_block_blocksize_1079 - 1)) begin
            write_burst_block_fsm_29 <= write_burst_block_fsm_29_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_1078 <= 1)) begin
            write_burst_block_fsm_29 <= write_burst_block_fsm_29_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_29 <= write_burst_block_fsm_29_init;
          end 
          if(0) begin
            write_burst_block_fsm_29 <= write_burst_block_fsm_29_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_30_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_30 <= write_burst_fsm_30_init;
      write_burst_addr_1086 <= 0;
      write_burst_stride_1087 <= 0;
      write_burst_length_1088 <= 0;
      write_burst_done_1089 <= 0;
    end else begin
      case(write_burst_fsm_30)
        write_burst_fsm_30_init: begin
          write_burst_addr_1086 <= _maxi_read_local_addr_buf;
          write_burst_stride_1087 <= _maxi_read_local_stride_buf;
          write_burst_length_1088 <= _maxi_read_local_size_buf;
          write_burst_done_1089 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 9) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_30 <= write_burst_fsm_30_1;
          end 
        end
        write_burst_fsm_30_1: begin
          if(write_burst_block_ram_wvalid_1084) begin
            write_burst_addr_1086 <= write_burst_addr_1086 + write_burst_stride_1087;
            write_burst_length_1088 <= write_burst_length_1088 - 1;
            write_burst_done_1089 <= 0;
          end 
          if(write_burst_block_ram_wvalid_1084 && (write_burst_length_1088 <= 1)) begin
            write_burst_done_1089 <= 1;
          end 
          if(write_burst_block_ram_wvalid_1084 && 0) begin
            write_burst_done_1089 <= 1;
          end 
          if(write_burst_block_ram_wvalid_1084 && (write_burst_length_1088 <= 1)) begin
            write_burst_fsm_30 <= write_burst_fsm_30_init;
          end 
          if(write_burst_block_ram_wvalid_1084 && 0) begin
            write_burst_fsm_30 <= write_burst_fsm_30_init;
          end 
          if(write_burst_block_ram_wquit_1085) begin
            write_burst_fsm_30 <= write_burst_fsm_30_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_31_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_31 <= write_burst_fsm_31_init;
      write_burst_addr_1092 <= 0;
      write_burst_stride_1093 <= 0;
      write_burst_length_1094 <= 0;
      write_burst_done_1095 <= 0;
    end else begin
      case(write_burst_fsm_31)
        write_burst_fsm_31_init: begin
          write_burst_addr_1092 <= _maxi_read_local_addr_buf;
          write_burst_stride_1093 <= _maxi_read_local_stride_buf;
          write_burst_length_1094 <= _maxi_read_local_size_buf;
          write_burst_done_1095 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 9) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_31 <= write_burst_fsm_31_1;
          end 
        end
        write_burst_fsm_31_1: begin
          if(write_burst_block_ram_wvalid_1090) begin
            write_burst_addr_1092 <= write_burst_addr_1092 + write_burst_stride_1093;
            write_burst_length_1094 <= write_burst_length_1094 - 1;
            write_burst_done_1095 <= 0;
          end 
          if(write_burst_block_ram_wvalid_1090 && (write_burst_length_1094 <= 1)) begin
            write_burst_done_1095 <= 1;
          end 
          if(write_burst_block_ram_wvalid_1090 && 0) begin
            write_burst_done_1095 <= 1;
          end 
          if(write_burst_block_ram_wvalid_1090 && (write_burst_length_1094 <= 1)) begin
            write_burst_fsm_31 <= write_burst_fsm_31_init;
          end 
          if(write_burst_block_ram_wvalid_1090 && 0) begin
            write_burst_fsm_31 <= write_burst_fsm_31_init;
          end 
          if(write_burst_block_ram_wquit_1091) begin
            write_burst_fsm_31 <= write_burst_fsm_31_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_32_1 = 1;
  localparam write_burst_block_fsm_32_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_32 <= write_burst_block_fsm_32_init;
      write_burst_block_length_1096 <= 0;
      write_burst_block_blocksize_1097 <= 0;
      write_burst_block_done_1098 <= 0;
      write_burst_block_count_1099 <= 0;
    end else begin
      case(write_burst_block_fsm_32)
        write_burst_block_fsm_32_init: begin
          write_burst_block_length_1096 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_1097 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_1098 <= 0;
          write_burst_block_count_1099 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 9) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_1;
          end 
        end
        write_burst_block_fsm_32_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_1096 <= write_burst_block_length_1096 - 1;
            write_burst_block_done_1098 <= 0;
            write_burst_block_count_1099 <= write_burst_block_count_1099 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_1096 <= 1)) begin
            write_burst_block_done_1098 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_1098 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_1099 == write_burst_block_blocksize_1097 - 1)) begin
            write_burst_block_count_1099 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_1099 == write_burst_block_blocksize_1097 - 1)) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_1096 <= 1)) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_init;
          end 
          if(0) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_init;
          end 
        end
        write_burst_block_fsm_32_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_1096 <= write_burst_block_length_1096 - 1;
            write_burst_block_done_1098 <= 0;
            write_burst_block_count_1099 <= write_burst_block_count_1099 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_1096 <= 1)) begin
            write_burst_block_done_1098 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_1098 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_1099 == write_burst_block_blocksize_1097 - 1)) begin
            write_burst_block_count_1099 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_1099 == write_burst_block_blocksize_1097 - 1)) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_1096 <= 1)) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_init;
          end 
          if(0) begin
            write_burst_block_fsm_32 <= write_burst_block_fsm_32_init;
          end 
        end
      endcase
    end
  end

  localparam max_pool_47_comp_fsm_1 = 1;
  localparam max_pool_47_comp_fsm_2 = 2;
  localparam max_pool_47_comp_fsm_3 = 3;
  localparam max_pool_47_comp_fsm_4 = 4;
  localparam max_pool_47_comp_fsm_5 = 5;
  localparam max_pool_47_comp_fsm_6 = 6;
  localparam max_pool_47_comp_fsm_7 = 7;

  always @(posedge CLK) begin
    if(RST) begin
      max_pool_47_comp_fsm <= max_pool_47_comp_fsm_init;
      max_pool_47_stream_act_local_0 <= 0;
      max_pool_47_stream_act_local_1 <= 0;
      max_pool_47_stream_act_local_2 <= 0;
      max_pool_47_stream_act_local_3 <= 0;
      max_pool_47_stream_out_local <= 0;
      max_pool_47_col_count <= 0;
      max_pool_47_col_select <= 0;
      max_pool_47_act_page_comp_offset_buf_0 <= 0;
      max_pool_47_act_page_comp_offset_buf_1 <= 0;
      max_pool_47_out_page_comp_offset_buf <= 0;
      max_pool_47_row_count_buf <= 0;
      max_pool_47_row_select_buf <= 0;
      max_pool_47_stream_pad_masks <= 0;
      max_pool_47_comp_count <= 0;
    end else begin
      if(control_max_pool_47 == 2) begin
        max_pool_47_comp_count <= 0;
      end 
      if(_stream_max_pool_47_sink_stop) begin
        max_pool_47_comp_count <= max_pool_47_comp_count + cparam_max_pool_47_inc_out_laddr;
      end 
      case(max_pool_47_comp_fsm)
        max_pool_47_comp_fsm_init: begin
          if((control_max_pool_47 == 12) && !max_pool_47_skip_comp) begin
            max_pool_47_comp_fsm <= max_pool_47_comp_fsm_1;
          end 
        end
        max_pool_47_comp_fsm_1: begin
          max_pool_47_stream_act_local_0 <= 0;
          if(cparam_max_pool_47_stream_act_local_small_flags_0) begin
            max_pool_47_stream_act_local_0 <= cparam_max_pool_47_stream_act_local_small_offset;
          end 
          if(cparam_max_pool_47_stream_act_local_large_flags_0) begin
            max_pool_47_stream_act_local_0 <= cparam_max_pool_47_stream_act_local_large_offset;
          end 
          max_pool_47_stream_act_local_1 <= 0;
          if(cparam_max_pool_47_stream_act_local_small_flags_1) begin
            max_pool_47_stream_act_local_1 <= cparam_max_pool_47_stream_act_local_small_offset;
          end 
          if(cparam_max_pool_47_stream_act_local_large_flags_1) begin
            max_pool_47_stream_act_local_1 <= cparam_max_pool_47_stream_act_local_large_offset;
          end 
          max_pool_47_stream_act_local_2 <= 0;
          if(cparam_max_pool_47_stream_act_local_small_flags_0) begin
            max_pool_47_stream_act_local_2 <= cparam_max_pool_47_stream_act_local_small_offset;
          end 
          if(cparam_max_pool_47_stream_act_local_large_flags_0) begin
            max_pool_47_stream_act_local_2 <= cparam_max_pool_47_stream_act_local_large_offset;
          end 
          max_pool_47_stream_act_local_3 <= 0;
          if(cparam_max_pool_47_stream_act_local_small_flags_1) begin
            max_pool_47_stream_act_local_3 <= cparam_max_pool_47_stream_act_local_small_offset;
          end 
          if(cparam_max_pool_47_stream_act_local_large_flags_1) begin
            max_pool_47_stream_act_local_3 <= cparam_max_pool_47_stream_act_local_large_offset;
          end 
          max_pool_47_stream_out_local <= 0;
          max_pool_47_col_count <= 0;
          max_pool_47_col_select <= cparam_max_pool_47_col_select_initval;
          max_pool_47_act_page_comp_offset_buf_0 <= max_pool_47_act_page_comp_offset_0;
          max_pool_47_act_page_comp_offset_buf_1 <= max_pool_47_act_page_comp_offset_1;
          max_pool_47_out_page_comp_offset_buf <= max_pool_47_out_page_comp_offset;
          max_pool_47_row_count_buf <= max_pool_47_row_count;
          max_pool_47_row_select_buf <= max_pool_47_row_select;
          max_pool_47_comp_fsm <= max_pool_47_comp_fsm_2;
        end
        max_pool_47_comp_fsm_2: begin
          max_pool_47_stream_pad_masks <= { (max_pool_47_row_select_buf == 0)? (max_pool_47_col_select == 0)? max_pool_47_stream_pad_mask_1_1 : 
                                          (max_pool_47_col_select == 1)? max_pool_47_stream_pad_mask_1_0 : 1'd0 : 
                                          (max_pool_47_row_select_buf == 1)? (max_pool_47_col_select == 0)? max_pool_47_stream_pad_mask_0_1 : 
                                          (max_pool_47_col_select == 1)? max_pool_47_stream_pad_mask_0_0 : 1'd0 : 1'd0, (max_pool_47_row_select_buf == 0)? (max_pool_47_col_select == 0)? max_pool_47_stream_pad_mask_1_0 : 
                                          (max_pool_47_col_select == 1)? max_pool_47_stream_pad_mask_1_1 : 1'd0 : 
                                          (max_pool_47_row_select_buf == 1)? (max_pool_47_col_select == 0)? max_pool_47_stream_pad_mask_0_0 : 
                                          (max_pool_47_col_select == 1)? max_pool_47_stream_pad_mask_0_1 : 1'd0 : 1'd0, (max_pool_47_row_select_buf == 0)? (max_pool_47_col_select == 0)? max_pool_47_stream_pad_mask_0_1 : 
                                          (max_pool_47_col_select == 1)? max_pool_47_stream_pad_mask_0_0 : 1'd0 : 
                                          (max_pool_47_row_select_buf == 1)? (max_pool_47_col_select == 0)? max_pool_47_stream_pad_mask_1_1 : 
                                          (max_pool_47_col_select == 1)? max_pool_47_stream_pad_mask_1_0 : 1'd0 : 1'd0, (max_pool_47_row_select_buf == 0)? (max_pool_47_col_select == 0)? max_pool_47_stream_pad_mask_0_0 : 
                                          (max_pool_47_col_select == 1)? max_pool_47_stream_pad_mask_0_1 : 1'd0 : 
                                          (max_pool_47_row_select_buf == 1)? (max_pool_47_col_select == 0)? max_pool_47_stream_pad_mask_1_0 : 
                                          (max_pool_47_col_select == 1)? max_pool_47_stream_pad_mask_1_1 : 1'd0 : 1'd0 };
          max_pool_47_comp_fsm <= max_pool_47_comp_fsm_3;
        end
        max_pool_47_comp_fsm_3: begin
          if(!_stream_max_pool_47_source_busy) begin
            max_pool_47_comp_fsm <= max_pool_47_comp_fsm_4;
          end 
        end
        max_pool_47_comp_fsm_4: begin
          max_pool_47_comp_fsm <= max_pool_47_comp_fsm_5;
          max_pool_47_comp_fsm <= max_pool_47_comp_fsm_5;
          max_pool_47_comp_fsm <= max_pool_47_comp_fsm_5;
          max_pool_47_comp_fsm <= max_pool_47_comp_fsm_5;
          max_pool_47_comp_fsm <= max_pool_47_comp_fsm_5;
          if(_stream_max_pool_47_stream_oready) begin
            max_pool_47_comp_fsm <= max_pool_47_comp_fsm_5;
          end 
        end
        max_pool_47_comp_fsm_5: begin
          max_pool_47_comp_fsm <= max_pool_47_comp_fsm_6;
        end
        max_pool_47_comp_fsm_6: begin
          if(_stream_max_pool_47_busy) begin
            max_pool_47_comp_fsm <= max_pool_47_comp_fsm_7;
          end 
        end
        max_pool_47_comp_fsm_7: begin
          if(!((max_pool_47_col_select == 0)? cparam_max_pool_47_inc_act_laddr_conds_0 : 
          (max_pool_47_col_select == 1)? cparam_max_pool_47_inc_act_laddr_conds_1 : 0)) begin
            max_pool_47_stream_act_local_0 <= max_pool_47_stream_act_local_0 + cparam_max_pool_47_inc_act_laddr_small;
          end 
          if((max_pool_47_col_select == 0)? cparam_max_pool_47_inc_act_laddr_conds_0 : 
          (max_pool_47_col_select == 1)? cparam_max_pool_47_inc_act_laddr_conds_1 : 0) begin
            max_pool_47_stream_act_local_0 <= max_pool_47_stream_act_local_0 + cparam_max_pool_47_inc_act_laddr_large;
          end 
          if(max_pool_47_col_count >= cparam_max_pool_47_max_col_count) begin
            max_pool_47_stream_act_local_0 <= 0;
          end 
          if((max_pool_47_col_count >= cparam_max_pool_47_max_col_count) && cparam_max_pool_47_stream_act_local_small_flags_0) begin
            max_pool_47_stream_act_local_0 <= cparam_max_pool_47_stream_act_local_small_offset;
          end 
          if((max_pool_47_col_count >= cparam_max_pool_47_max_col_count) && cparam_max_pool_47_stream_act_local_large_flags_0) begin
            max_pool_47_stream_act_local_0 <= cparam_max_pool_47_stream_act_local_large_offset;
          end 
          if(!((max_pool_47_col_select == 0)? cparam_max_pool_47_inc_act_laddr_conds_2 : 
          (max_pool_47_col_select == 1)? cparam_max_pool_47_inc_act_laddr_conds_3 : 0)) begin
            max_pool_47_stream_act_local_1 <= max_pool_47_stream_act_local_1 + cparam_max_pool_47_inc_act_laddr_small;
          end 
          if((max_pool_47_col_select == 0)? cparam_max_pool_47_inc_act_laddr_conds_2 : 
          (max_pool_47_col_select == 1)? cparam_max_pool_47_inc_act_laddr_conds_3 : 0) begin
            max_pool_47_stream_act_local_1 <= max_pool_47_stream_act_local_1 + cparam_max_pool_47_inc_act_laddr_large;
          end 
          if(max_pool_47_col_count >= cparam_max_pool_47_max_col_count) begin
            max_pool_47_stream_act_local_1 <= 0;
          end 
          if((max_pool_47_col_count >= cparam_max_pool_47_max_col_count) && cparam_max_pool_47_stream_act_local_small_flags_1) begin
            max_pool_47_stream_act_local_1 <= cparam_max_pool_47_stream_act_local_small_offset;
          end 
          if((max_pool_47_col_count >= cparam_max_pool_47_max_col_count) && cparam_max_pool_47_stream_act_local_large_flags_1) begin
            max_pool_47_stream_act_local_1 <= cparam_max_pool_47_stream_act_local_large_offset;
          end 
          if(!((max_pool_47_col_select == 0)? cparam_max_pool_47_inc_act_laddr_conds_4 : 
          (max_pool_47_col_select == 1)? cparam_max_pool_47_inc_act_laddr_conds_5 : 0)) begin
            max_pool_47_stream_act_local_2 <= max_pool_47_stream_act_local_2 + cparam_max_pool_47_inc_act_laddr_small;
          end 
          if((max_pool_47_col_select == 0)? cparam_max_pool_47_inc_act_laddr_conds_4 : 
          (max_pool_47_col_select == 1)? cparam_max_pool_47_inc_act_laddr_conds_5 : 0) begin
            max_pool_47_stream_act_local_2 <= max_pool_47_stream_act_local_2 + cparam_max_pool_47_inc_act_laddr_large;
          end 
          if(max_pool_47_col_count >= cparam_max_pool_47_max_col_count) begin
            max_pool_47_stream_act_local_2 <= 0;
          end 
          if((max_pool_47_col_count >= cparam_max_pool_47_max_col_count) && cparam_max_pool_47_stream_act_local_small_flags_0) begin
            max_pool_47_stream_act_local_2 <= cparam_max_pool_47_stream_act_local_small_offset;
          end 
          if((max_pool_47_col_count >= cparam_max_pool_47_max_col_count) && cparam_max_pool_47_stream_act_local_large_flags_0) begin
            max_pool_47_stream_act_local_2 <= cparam_max_pool_47_stream_act_local_large_offset;
          end 
          if(!((max_pool_47_col_select == 0)? cparam_max_pool_47_inc_act_laddr_conds_6 : 
          (max_pool_47_col_select == 1)? cparam_max_pool_47_inc_act_laddr_conds_7 : 0)) begin
            max_pool_47_stream_act_local_3 <= max_pool_47_stream_act_local_3 + cparam_max_pool_47_inc_act_laddr_small;
          end 
          if((max_pool_47_col_select == 0)? cparam_max_pool_47_inc_act_laddr_conds_6 : 
          (max_pool_47_col_select == 1)? cparam_max_pool_47_inc_act_laddr_conds_7 : 0) begin
            max_pool_47_stream_act_local_3 <= max_pool_47_stream_act_local_3 + cparam_max_pool_47_inc_act_laddr_large;
          end 
          if(max_pool_47_col_count >= cparam_max_pool_47_max_col_count) begin
            max_pool_47_stream_act_local_3 <= 0;
          end 
          if((max_pool_47_col_count >= cparam_max_pool_47_max_col_count) && cparam_max_pool_47_stream_act_local_small_flags_1) begin
            max_pool_47_stream_act_local_3 <= cparam_max_pool_47_stream_act_local_small_offset;
          end 
          if((max_pool_47_col_count >= cparam_max_pool_47_max_col_count) && cparam_max_pool_47_stream_act_local_large_flags_1) begin
            max_pool_47_stream_act_local_3 <= cparam_max_pool_47_stream_act_local_large_offset;
          end 
          max_pool_47_stream_out_local <= max_pool_47_stream_out_local + cparam_max_pool_47_inc_out_laddr;
          if(max_pool_47_col_count >= cparam_max_pool_47_max_col_count) begin
            max_pool_47_stream_out_local <= 0;
          end 
          max_pool_47_col_count <= max_pool_47_col_count + cparam_max_pool_47_stride_col;
          if(max_pool_47_col_count >= cparam_max_pool_47_max_col_count) begin
            max_pool_47_col_count <= 0;
          end 
          max_pool_47_col_select <= max_pool_47_col_select + cparam_max_pool_47_stride_col_mod_ksize;
          if(max_pool_47_col_select + cparam_max_pool_47_stride_col_mod_ksize >= 2) begin
            max_pool_47_col_select <= max_pool_47_col_select - cparam_max_pool_47_ksize_col_minus_stride_col_mod;
          end 
          if(max_pool_47_col_count >= cparam_max_pool_47_max_col_count) begin
            max_pool_47_col_select <= cparam_max_pool_47_col_select_initval;
          end 
          max_pool_47_comp_fsm <= max_pool_47_comp_fsm_2;
          if(max_pool_47_col_count >= cparam_max_pool_47_max_col_count) begin
            max_pool_47_comp_fsm <= max_pool_47_comp_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_max_pool_47_source_1_source_fsm_0_1 = 1;
  localparam _stream_max_pool_47_source_1_source_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_47_source_1_source_fsm_0 <= _stream_max_pool_47_source_1_source_fsm_0_init;
    end else begin
      case(_stream_max_pool_47_source_1_source_fsm_0)
        _stream_max_pool_47_source_1_source_fsm_0_init: begin
          if(_stream_max_pool_47_source_start && _stream_max_pool_47_source_1_source_mode & 5'b1 && _stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_source_1_source_fsm_0 <= _stream_max_pool_47_source_1_source_fsm_0_1;
          end 
        end
        _stream_max_pool_47_source_1_source_fsm_0_1: begin
          if(_stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_source_1_source_fsm_0 <= _stream_max_pool_47_source_1_source_fsm_0_2;
          end 
        end
        _stream_max_pool_47_source_1_source_fsm_0_2: begin
          if((_stream_max_pool_47_source_1_source_count == 1) && _stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_source_1_source_fsm_0 <= _stream_max_pool_47_source_1_source_fsm_0_init;
          end 
          if(_stream_max_pool_47_source_stop && _stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_source_1_source_fsm_0 <= _stream_max_pool_47_source_1_source_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_max_pool_47_source_2_source_fsm_1_1 = 1;
  localparam _stream_max_pool_47_source_2_source_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_47_source_2_source_fsm_1 <= _stream_max_pool_47_source_2_source_fsm_1_init;
    end else begin
      case(_stream_max_pool_47_source_2_source_fsm_1)
        _stream_max_pool_47_source_2_source_fsm_1_init: begin
          if(_stream_max_pool_47_source_start && _stream_max_pool_47_source_2_source_mode & 5'b1 && _stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_source_2_source_fsm_1 <= _stream_max_pool_47_source_2_source_fsm_1_1;
          end 
        end
        _stream_max_pool_47_source_2_source_fsm_1_1: begin
          if(_stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_source_2_source_fsm_1 <= _stream_max_pool_47_source_2_source_fsm_1_2;
          end 
        end
        _stream_max_pool_47_source_2_source_fsm_1_2: begin
          if((_stream_max_pool_47_source_2_source_count == 1) && _stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_source_2_source_fsm_1 <= _stream_max_pool_47_source_2_source_fsm_1_init;
          end 
          if(_stream_max_pool_47_source_stop && _stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_source_2_source_fsm_1 <= _stream_max_pool_47_source_2_source_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_max_pool_47_source_3_source_fsm_2_1 = 1;
  localparam _stream_max_pool_47_source_3_source_fsm_2_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_47_source_3_source_fsm_2 <= _stream_max_pool_47_source_3_source_fsm_2_init;
    end else begin
      case(_stream_max_pool_47_source_3_source_fsm_2)
        _stream_max_pool_47_source_3_source_fsm_2_init: begin
          if(_stream_max_pool_47_source_start && _stream_max_pool_47_source_3_source_mode & 5'b1 && _stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_source_3_source_fsm_2 <= _stream_max_pool_47_source_3_source_fsm_2_1;
          end 
        end
        _stream_max_pool_47_source_3_source_fsm_2_1: begin
          if(_stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_source_3_source_fsm_2 <= _stream_max_pool_47_source_3_source_fsm_2_2;
          end 
        end
        _stream_max_pool_47_source_3_source_fsm_2_2: begin
          if((_stream_max_pool_47_source_3_source_count == 1) && _stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_source_3_source_fsm_2 <= _stream_max_pool_47_source_3_source_fsm_2_init;
          end 
          if(_stream_max_pool_47_source_stop && _stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_source_3_source_fsm_2 <= _stream_max_pool_47_source_3_source_fsm_2_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_max_pool_47_source_4_source_fsm_3_1 = 1;
  localparam _stream_max_pool_47_source_4_source_fsm_3_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_47_source_4_source_fsm_3 <= _stream_max_pool_47_source_4_source_fsm_3_init;
    end else begin
      case(_stream_max_pool_47_source_4_source_fsm_3)
        _stream_max_pool_47_source_4_source_fsm_3_init: begin
          if(_stream_max_pool_47_source_start && _stream_max_pool_47_source_4_source_mode & 5'b1 && _stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_source_4_source_fsm_3 <= _stream_max_pool_47_source_4_source_fsm_3_1;
          end 
        end
        _stream_max_pool_47_source_4_source_fsm_3_1: begin
          if(_stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_source_4_source_fsm_3 <= _stream_max_pool_47_source_4_source_fsm_3_2;
          end 
        end
        _stream_max_pool_47_source_4_source_fsm_3_2: begin
          if((_stream_max_pool_47_source_4_source_count == 1) && _stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_source_4_source_fsm_3 <= _stream_max_pool_47_source_4_source_fsm_3_init;
          end 
          if(_stream_max_pool_47_source_stop && _stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_source_4_source_fsm_3 <= _stream_max_pool_47_source_4_source_fsm_3_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_max_pool_47_sink_6_sink_fsm_4_1 = 1;
  localparam _stream_max_pool_47_sink_6_sink_fsm_4_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_47_sink_6_sink_fsm_4 <= _stream_max_pool_47_sink_6_sink_fsm_4_init;
    end else begin
      case(_stream_max_pool_47_sink_6_sink_fsm_4)
        _stream_max_pool_47_sink_6_sink_fsm_4_init: begin
          if(_stream_max_pool_47_sink_start && _stream_max_pool_47_sink_6_sink_mode & 5'b1 && _stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_sink_6_sink_fsm_4 <= _stream_max_pool_47_sink_6_sink_fsm_4_1;
          end 
        end
        _stream_max_pool_47_sink_6_sink_fsm_4_1: begin
          if(_stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_sink_6_sink_fsm_4 <= _stream_max_pool_47_sink_6_sink_fsm_4_2;
          end 
        end
        _stream_max_pool_47_sink_6_sink_fsm_4_2: begin
          if((_stream_max_pool_47_sink_6_sink_count == 1) && _stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_sink_6_sink_fsm_4 <= _stream_max_pool_47_sink_6_sink_fsm_4_init;
          end 
          if(_stream_max_pool_47_sink_stop && _stream_max_pool_47_stream_oready) begin
            _stream_max_pool_47_sink_6_sink_fsm_4 <= _stream_max_pool_47_sink_6_sink_fsm_4_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_fsm_33_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_fsm_33 <= read_burst_fsm_33_init;
      read_burst_addr_1196 <= 0;
      read_burst_stride_1197 <= 0;
      read_burst_length_1198 <= 0;
      read_burst_rvalid_1199 <= 0;
      read_burst_rlast_1200 <= 0;
    end else begin
      case(read_burst_fsm_33)
        read_burst_fsm_33_init: begin
          read_burst_addr_1196 <= _maxi_write_local_addr_buf;
          read_burst_stride_1197 <= _maxi_write_local_stride_buf;
          read_burst_length_1198 <= _maxi_write_size_buf;
          read_burst_rvalid_1199 <= 0;
          read_burst_rlast_1200 <= 0;
          if((_maxi_write_data_fsm == 1) && (_maxi_write_op_sel_buf == 3) && (_maxi_write_size_buf > 0)) begin
            read_burst_fsm_33 <= read_burst_fsm_33_1;
          end 
        end
        read_burst_fsm_33_1: begin
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_length_1198 > 0)) begin
            read_burst_addr_1196 <= read_burst_addr_1196 + read_burst_stride_1197;
            read_burst_length_1198 <= read_burst_length_1198 - 1;
            read_burst_rvalid_1199 <= 1;
          end 
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_length_1198 <= 1)) begin
            read_burst_rlast_1200 <= 1;
          end 
          if(read_burst_rlast_1200 && read_burst_rvalid_1199 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_rvalid_1199 <= 0;
            read_burst_rlast_1200 <= 0;
          end 
          if(0) begin
            read_burst_rvalid_1199 <= 0;
            read_burst_rlast_1200 <= 0;
          end 
          if(read_burst_rlast_1200 && read_burst_rvalid_1199 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_fsm_33 <= read_burst_fsm_33_init;
          end 
          if(0) begin
            read_burst_fsm_33 <= read_burst_fsm_33_init;
          end 
        end
      endcase
    end
  end


endmodule



module _maxi_read_req_fifo
(
  input CLK,
  input RST,
  input _maxi_read_req_fifo_enq,
  input [137-1:0] _maxi_read_req_fifo_wdata,
  output _maxi_read_req_fifo_full,
  output _maxi_read_req_fifo_almost_full,
  input _maxi_read_req_fifo_deq,
  output [137-1:0] _maxi_read_req_fifo_rdata,
  output _maxi_read_req_fifo_empty,
  output _maxi_read_req_fifo_almost_empty
);

  reg [137-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [137-1:0] rdata;
  assign _maxi_read_req_fifo_full = is_full;
  assign _maxi_read_req_fifo_almost_full = is_almost_full || is_full;
  assign _maxi_read_req_fifo_empty = is_empty;
  assign _maxi_read_req_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _maxi_read_req_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_maxi_read_req_fifo_enq && !is_full) begin
        mem[head] <= _maxi_read_req_fifo_wdata;
        head <= head + 1;
      end 
      if(_maxi_read_req_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module _maxi_write_req_fifo
(
  input CLK,
  input RST,
  input _maxi_write_req_fifo_enq,
  input [137-1:0] _maxi_write_req_fifo_wdata,
  output _maxi_write_req_fifo_full,
  output _maxi_write_req_fifo_almost_full,
  input _maxi_write_req_fifo_deq,
  output [137-1:0] _maxi_write_req_fifo_rdata,
  output _maxi_write_req_fifo_empty,
  output _maxi_write_req_fifo_almost_empty
);

  reg [137-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [137-1:0] rdata;
  assign _maxi_write_req_fifo_full = is_full;
  assign _maxi_write_req_fifo_almost_full = is_almost_full || is_full;
  assign _maxi_write_req_fifo_empty = is_empty;
  assign _maxi_write_req_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _maxi_write_req_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_maxi_write_req_fifo_enq && !is_full) begin
        mem[head] <= _maxi_write_req_fifo_wdata;
        head <= head + 1;
      end 
      if(_maxi_write_req_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module ram_w32_l32768_id0
(
  input CLK,
  input [15-1:0] ram_w32_l32768_id0_0_addr,
  output [32-1:0] ram_w32_l32768_id0_0_rdata,
  input [32-1:0] ram_w32_l32768_id0_0_wdata,
  input ram_w32_l32768_id0_0_wenable,
  input ram_w32_l32768_id0_0_enable,
  input [15-1:0] ram_w32_l32768_id0_1_addr,
  output [32-1:0] ram_w32_l32768_id0_1_rdata,
  input [32-1:0] ram_w32_l32768_id0_1_wdata,
  input ram_w32_l32768_id0_1_wenable,
  input ram_w32_l32768_id0_1_enable
);

  reg [32-1:0] ram_w32_l32768_id0_0_rdata_out;
  assign ram_w32_l32768_id0_0_rdata = ram_w32_l32768_id0_0_rdata_out;
  reg [32-1:0] ram_w32_l32768_id0_1_rdata_out;
  assign ram_w32_l32768_id0_1_rdata = ram_w32_l32768_id0_1_rdata_out;
  reg [32-1:0] mem [0:32768-1];

  always @(posedge CLK) begin
    if(ram_w32_l32768_id0_0_enable) begin
      if(ram_w32_l32768_id0_0_wenable) begin
        mem[ram_w32_l32768_id0_0_addr] <= ram_w32_l32768_id0_0_wdata;
        ram_w32_l32768_id0_0_rdata_out <= ram_w32_l32768_id0_0_wdata;
      end else begin
        ram_w32_l32768_id0_0_rdata_out <= mem[ram_w32_l32768_id0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l32768_id0_1_enable) begin
      if(ram_w32_l32768_id0_1_wenable) begin
        mem[ram_w32_l32768_id0_1_addr] <= ram_w32_l32768_id0_1_wdata;
        ram_w32_l32768_id0_1_rdata_out <= ram_w32_l32768_id0_1_wdata;
      end else begin
        ram_w32_l32768_id0_1_rdata_out <= mem[ram_w32_l32768_id0_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l16384_id0
(
  input CLK,
  input [14-1:0] ram_w32_l16384_id0_0_addr,
  output [32-1:0] ram_w32_l16384_id0_0_rdata,
  input [32-1:0] ram_w32_l16384_id0_0_wdata,
  input ram_w32_l16384_id0_0_wenable,
  input ram_w32_l16384_id0_0_enable,
  input [14-1:0] ram_w32_l16384_id0_1_addr,
  output [32-1:0] ram_w32_l16384_id0_1_rdata,
  input [32-1:0] ram_w32_l16384_id0_1_wdata,
  input ram_w32_l16384_id0_1_wenable,
  input ram_w32_l16384_id0_1_enable
);

  reg [32-1:0] ram_w32_l16384_id0_0_rdata_out;
  assign ram_w32_l16384_id0_0_rdata = ram_w32_l16384_id0_0_rdata_out;
  reg [32-1:0] ram_w32_l16384_id0_1_rdata_out;
  assign ram_w32_l16384_id0_1_rdata = ram_w32_l16384_id0_1_rdata_out;
  reg [32-1:0] mem [0:16384-1];

  always @(posedge CLK) begin
    if(ram_w32_l16384_id0_0_enable) begin
      if(ram_w32_l16384_id0_0_wenable) begin
        mem[ram_w32_l16384_id0_0_addr] <= ram_w32_l16384_id0_0_wdata;
        ram_w32_l16384_id0_0_rdata_out <= ram_w32_l16384_id0_0_wdata;
      end else begin
        ram_w32_l16384_id0_0_rdata_out <= mem[ram_w32_l16384_id0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l16384_id0_1_enable) begin
      if(ram_w32_l16384_id0_1_wenable) begin
        mem[ram_w32_l16384_id0_1_addr] <= ram_w32_l16384_id0_1_wdata;
        ram_w32_l16384_id0_1_rdata_out <= ram_w32_l16384_id0_1_wdata;
      end else begin
        ram_w32_l16384_id0_1_rdata_out <= mem[ram_w32_l16384_id0_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l8192_id0
(
  input CLK,
  input [13-1:0] ram_w32_l8192_id0_0_addr,
  output [32-1:0] ram_w32_l8192_id0_0_rdata,
  input [32-1:0] ram_w32_l8192_id0_0_wdata,
  input ram_w32_l8192_id0_0_wenable,
  input ram_w32_l8192_id0_0_enable,
  input [13-1:0] ram_w32_l8192_id0_1_addr,
  output [32-1:0] ram_w32_l8192_id0_1_rdata,
  input [32-1:0] ram_w32_l8192_id0_1_wdata,
  input ram_w32_l8192_id0_1_wenable,
  input ram_w32_l8192_id0_1_enable
);

  reg [32-1:0] ram_w32_l8192_id0_0_rdata_out;
  assign ram_w32_l8192_id0_0_rdata = ram_w32_l8192_id0_0_rdata_out;
  reg [32-1:0] ram_w32_l8192_id0_1_rdata_out;
  assign ram_w32_l8192_id0_1_rdata = ram_w32_l8192_id0_1_rdata_out;
  reg [32-1:0] mem [0:8192-1];

  always @(posedge CLK) begin
    if(ram_w32_l8192_id0_0_enable) begin
      if(ram_w32_l8192_id0_0_wenable) begin
        mem[ram_w32_l8192_id0_0_addr] <= ram_w32_l8192_id0_0_wdata;
        ram_w32_l8192_id0_0_rdata_out <= ram_w32_l8192_id0_0_wdata;
      end else begin
        ram_w32_l8192_id0_0_rdata_out <= mem[ram_w32_l8192_id0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l8192_id0_1_enable) begin
      if(ram_w32_l8192_id0_1_wenable) begin
        mem[ram_w32_l8192_id0_1_addr] <= ram_w32_l8192_id0_1_wdata;
        ram_w32_l8192_id0_1_rdata_out <= ram_w32_l8192_id0_1_wdata;
      end else begin
        ram_w32_l8192_id0_1_rdata_out <= mem[ram_w32_l8192_id0_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l8192_id1
(
  input CLK,
  input [13-1:0] ram_w32_l8192_id1_0_addr,
  output [32-1:0] ram_w32_l8192_id1_0_rdata,
  input [32-1:0] ram_w32_l8192_id1_0_wdata,
  input ram_w32_l8192_id1_0_wenable,
  input ram_w32_l8192_id1_0_enable,
  input [13-1:0] ram_w32_l8192_id1_1_addr,
  output [32-1:0] ram_w32_l8192_id1_1_rdata,
  input [32-1:0] ram_w32_l8192_id1_1_wdata,
  input ram_w32_l8192_id1_1_wenable,
  input ram_w32_l8192_id1_1_enable
);

  reg [32-1:0] ram_w32_l8192_id1_0_rdata_out;
  assign ram_w32_l8192_id1_0_rdata = ram_w32_l8192_id1_0_rdata_out;
  reg [32-1:0] ram_w32_l8192_id1_1_rdata_out;
  assign ram_w32_l8192_id1_1_rdata = ram_w32_l8192_id1_1_rdata_out;
  reg [32-1:0] mem [0:8192-1];

  always @(posedge CLK) begin
    if(ram_w32_l8192_id1_0_enable) begin
      if(ram_w32_l8192_id1_0_wenable) begin
        mem[ram_w32_l8192_id1_0_addr] <= ram_w32_l8192_id1_0_wdata;
        ram_w32_l8192_id1_0_rdata_out <= ram_w32_l8192_id1_0_wdata;
      end else begin
        ram_w32_l8192_id1_0_rdata_out <= mem[ram_w32_l8192_id1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l8192_id1_1_enable) begin
      if(ram_w32_l8192_id1_1_wenable) begin
        mem[ram_w32_l8192_id1_1_addr] <= ram_w32_l8192_id1_1_wdata;
        ram_w32_l8192_id1_1_rdata_out <= ram_w32_l8192_id1_1_wdata;
      end else begin
        ram_w32_l8192_id1_1_rdata_out <= mem[ram_w32_l8192_id1_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l8192_id2
(
  input CLK,
  input [13-1:0] ram_w32_l8192_id2_0_addr,
  output [32-1:0] ram_w32_l8192_id2_0_rdata,
  input [32-1:0] ram_w32_l8192_id2_0_wdata,
  input ram_w32_l8192_id2_0_wenable,
  input ram_w32_l8192_id2_0_enable,
  input [13-1:0] ram_w32_l8192_id2_1_addr,
  output [32-1:0] ram_w32_l8192_id2_1_rdata,
  input [32-1:0] ram_w32_l8192_id2_1_wdata,
  input ram_w32_l8192_id2_1_wenable,
  input ram_w32_l8192_id2_1_enable
);

  reg [32-1:0] ram_w32_l8192_id2_0_rdata_out;
  assign ram_w32_l8192_id2_0_rdata = ram_w32_l8192_id2_0_rdata_out;
  reg [32-1:0] ram_w32_l8192_id2_1_rdata_out;
  assign ram_w32_l8192_id2_1_rdata = ram_w32_l8192_id2_1_rdata_out;
  reg [32-1:0] mem [0:8192-1];

  always @(posedge CLK) begin
    if(ram_w32_l8192_id2_0_enable) begin
      if(ram_w32_l8192_id2_0_wenable) begin
        mem[ram_w32_l8192_id2_0_addr] <= ram_w32_l8192_id2_0_wdata;
        ram_w32_l8192_id2_0_rdata_out <= ram_w32_l8192_id2_0_wdata;
      end else begin
        ram_w32_l8192_id2_0_rdata_out <= mem[ram_w32_l8192_id2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l8192_id2_1_enable) begin
      if(ram_w32_l8192_id2_1_wenable) begin
        mem[ram_w32_l8192_id2_1_addr] <= ram_w32_l8192_id2_1_wdata;
        ram_w32_l8192_id2_1_rdata_out <= ram_w32_l8192_id2_1_wdata;
      end else begin
        ram_w32_l8192_id2_1_rdata_out <= mem[ram_w32_l8192_id2_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l8192_id3
(
  input CLK,
  input [13-1:0] ram_w32_l8192_id3_0_addr,
  output [32-1:0] ram_w32_l8192_id3_0_rdata,
  input [32-1:0] ram_w32_l8192_id3_0_wdata,
  input ram_w32_l8192_id3_0_wenable,
  input ram_w32_l8192_id3_0_enable,
  input [13-1:0] ram_w32_l8192_id3_1_addr,
  output [32-1:0] ram_w32_l8192_id3_1_rdata,
  input [32-1:0] ram_w32_l8192_id3_1_wdata,
  input ram_w32_l8192_id3_1_wenable,
  input ram_w32_l8192_id3_1_enable
);

  reg [32-1:0] ram_w32_l8192_id3_0_rdata_out;
  assign ram_w32_l8192_id3_0_rdata = ram_w32_l8192_id3_0_rdata_out;
  reg [32-1:0] ram_w32_l8192_id3_1_rdata_out;
  assign ram_w32_l8192_id3_1_rdata = ram_w32_l8192_id3_1_rdata_out;
  reg [32-1:0] mem [0:8192-1];

  always @(posedge CLK) begin
    if(ram_w32_l8192_id3_0_enable) begin
      if(ram_w32_l8192_id3_0_wenable) begin
        mem[ram_w32_l8192_id3_0_addr] <= ram_w32_l8192_id3_0_wdata;
        ram_w32_l8192_id3_0_rdata_out <= ram_w32_l8192_id3_0_wdata;
      end else begin
        ram_w32_l8192_id3_0_rdata_out <= mem[ram_w32_l8192_id3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l8192_id3_1_enable) begin
      if(ram_w32_l8192_id3_1_wenable) begin
        mem[ram_w32_l8192_id3_1_addr] <= ram_w32_l8192_id3_1_wdata;
        ram_w32_l8192_id3_1_rdata_out <= ram_w32_l8192_id3_1_wdata;
      end else begin
        ram_w32_l8192_id3_1_rdata_out <= mem[ram_w32_l8192_id3_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l4096_id0
(
  input CLK,
  input [12-1:0] ram_w32_l4096_id0_0_addr,
  output [32-1:0] ram_w32_l4096_id0_0_rdata,
  input [32-1:0] ram_w32_l4096_id0_0_wdata,
  input ram_w32_l4096_id0_0_wenable,
  input ram_w32_l4096_id0_0_enable,
  input [12-1:0] ram_w32_l4096_id0_1_addr,
  output [32-1:0] ram_w32_l4096_id0_1_rdata,
  input [32-1:0] ram_w32_l4096_id0_1_wdata,
  input ram_w32_l4096_id0_1_wenable,
  input ram_w32_l4096_id0_1_enable
);

  reg [32-1:0] ram_w32_l4096_id0_0_rdata_out;
  assign ram_w32_l4096_id0_0_rdata = ram_w32_l4096_id0_0_rdata_out;
  reg [32-1:0] ram_w32_l4096_id0_1_rdata_out;
  assign ram_w32_l4096_id0_1_rdata = ram_w32_l4096_id0_1_rdata_out;
  reg [32-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w32_l4096_id0_0_enable) begin
      if(ram_w32_l4096_id0_0_wenable) begin
        mem[ram_w32_l4096_id0_0_addr] <= ram_w32_l4096_id0_0_wdata;
        ram_w32_l4096_id0_0_rdata_out <= ram_w32_l4096_id0_0_wdata;
      end else begin
        ram_w32_l4096_id0_0_rdata_out <= mem[ram_w32_l4096_id0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l4096_id0_1_enable) begin
      if(ram_w32_l4096_id0_1_wenable) begin
        mem[ram_w32_l4096_id0_1_addr] <= ram_w32_l4096_id0_1_wdata;
        ram_w32_l4096_id0_1_rdata_out <= ram_w32_l4096_id0_1_wdata;
      end else begin
        ram_w32_l4096_id0_1_rdata_out <= mem[ram_w32_l4096_id0_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l4096_id1
(
  input CLK,
  input [12-1:0] ram_w32_l4096_id1_0_addr,
  output [32-1:0] ram_w32_l4096_id1_0_rdata,
  input [32-1:0] ram_w32_l4096_id1_0_wdata,
  input ram_w32_l4096_id1_0_wenable,
  input ram_w32_l4096_id1_0_enable,
  input [12-1:0] ram_w32_l4096_id1_1_addr,
  output [32-1:0] ram_w32_l4096_id1_1_rdata,
  input [32-1:0] ram_w32_l4096_id1_1_wdata,
  input ram_w32_l4096_id1_1_wenable,
  input ram_w32_l4096_id1_1_enable
);

  reg [32-1:0] ram_w32_l4096_id1_0_rdata_out;
  assign ram_w32_l4096_id1_0_rdata = ram_w32_l4096_id1_0_rdata_out;
  reg [32-1:0] ram_w32_l4096_id1_1_rdata_out;
  assign ram_w32_l4096_id1_1_rdata = ram_w32_l4096_id1_1_rdata_out;
  reg [32-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w32_l4096_id1_0_enable) begin
      if(ram_w32_l4096_id1_0_wenable) begin
        mem[ram_w32_l4096_id1_0_addr] <= ram_w32_l4096_id1_0_wdata;
        ram_w32_l4096_id1_0_rdata_out <= ram_w32_l4096_id1_0_wdata;
      end else begin
        ram_w32_l4096_id1_0_rdata_out <= mem[ram_w32_l4096_id1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l4096_id1_1_enable) begin
      if(ram_w32_l4096_id1_1_wenable) begin
        mem[ram_w32_l4096_id1_1_addr] <= ram_w32_l4096_id1_1_wdata;
        ram_w32_l4096_id1_1_rdata_out <= ram_w32_l4096_id1_1_wdata;
      end else begin
        ram_w32_l4096_id1_1_rdata_out <= mem[ram_w32_l4096_id1_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l4096_id2
(
  input CLK,
  input [12-1:0] ram_w32_l4096_id2_0_addr,
  output [32-1:0] ram_w32_l4096_id2_0_rdata,
  input [32-1:0] ram_w32_l4096_id2_0_wdata,
  input ram_w32_l4096_id2_0_wenable,
  input ram_w32_l4096_id2_0_enable,
  input [12-1:0] ram_w32_l4096_id2_1_addr,
  output [32-1:0] ram_w32_l4096_id2_1_rdata,
  input [32-1:0] ram_w32_l4096_id2_1_wdata,
  input ram_w32_l4096_id2_1_wenable,
  input ram_w32_l4096_id2_1_enable
);

  reg [32-1:0] ram_w32_l4096_id2_0_rdata_out;
  assign ram_w32_l4096_id2_0_rdata = ram_w32_l4096_id2_0_rdata_out;
  reg [32-1:0] ram_w32_l4096_id2_1_rdata_out;
  assign ram_w32_l4096_id2_1_rdata = ram_w32_l4096_id2_1_rdata_out;
  reg [32-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w32_l4096_id2_0_enable) begin
      if(ram_w32_l4096_id2_0_wenable) begin
        mem[ram_w32_l4096_id2_0_addr] <= ram_w32_l4096_id2_0_wdata;
        ram_w32_l4096_id2_0_rdata_out <= ram_w32_l4096_id2_0_wdata;
      end else begin
        ram_w32_l4096_id2_0_rdata_out <= mem[ram_w32_l4096_id2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l4096_id2_1_enable) begin
      if(ram_w32_l4096_id2_1_wenable) begin
        mem[ram_w32_l4096_id2_1_addr] <= ram_w32_l4096_id2_1_wdata;
        ram_w32_l4096_id2_1_rdata_out <= ram_w32_l4096_id2_1_wdata;
      end else begin
        ram_w32_l4096_id2_1_rdata_out <= mem[ram_w32_l4096_id2_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l4096_id3
(
  input CLK,
  input [12-1:0] ram_w32_l4096_id3_0_addr,
  output [32-1:0] ram_w32_l4096_id3_0_rdata,
  input [32-1:0] ram_w32_l4096_id3_0_wdata,
  input ram_w32_l4096_id3_0_wenable,
  input ram_w32_l4096_id3_0_enable,
  input [12-1:0] ram_w32_l4096_id3_1_addr,
  output [32-1:0] ram_w32_l4096_id3_1_rdata,
  input [32-1:0] ram_w32_l4096_id3_1_wdata,
  input ram_w32_l4096_id3_1_wenable,
  input ram_w32_l4096_id3_1_enable
);

  reg [32-1:0] ram_w32_l4096_id3_0_rdata_out;
  assign ram_w32_l4096_id3_0_rdata = ram_w32_l4096_id3_0_rdata_out;
  reg [32-1:0] ram_w32_l4096_id3_1_rdata_out;
  assign ram_w32_l4096_id3_1_rdata = ram_w32_l4096_id3_1_rdata_out;
  reg [32-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w32_l4096_id3_0_enable) begin
      if(ram_w32_l4096_id3_0_wenable) begin
        mem[ram_w32_l4096_id3_0_addr] <= ram_w32_l4096_id3_0_wdata;
        ram_w32_l4096_id3_0_rdata_out <= ram_w32_l4096_id3_0_wdata;
      end else begin
        ram_w32_l4096_id3_0_rdata_out <= mem[ram_w32_l4096_id3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l4096_id3_1_enable) begin
      if(ram_w32_l4096_id3_1_wenable) begin
        mem[ram_w32_l4096_id3_1_addr] <= ram_w32_l4096_id3_1_wdata;
        ram_w32_l4096_id3_1_rdata_out <= ram_w32_l4096_id3_1_wdata;
      end else begin
        ram_w32_l4096_id3_1_rdata_out <= mem[ram_w32_l4096_id3_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l4096_id4
(
  input CLK,
  input [12-1:0] ram_w32_l4096_id4_0_addr,
  output [32-1:0] ram_w32_l4096_id4_0_rdata,
  input [32-1:0] ram_w32_l4096_id4_0_wdata,
  input ram_w32_l4096_id4_0_wenable,
  input ram_w32_l4096_id4_0_enable,
  input [12-1:0] ram_w32_l4096_id4_1_addr,
  output [32-1:0] ram_w32_l4096_id4_1_rdata,
  input [32-1:0] ram_w32_l4096_id4_1_wdata,
  input ram_w32_l4096_id4_1_wenable,
  input ram_w32_l4096_id4_1_enable
);

  reg [32-1:0] ram_w32_l4096_id4_0_rdata_out;
  assign ram_w32_l4096_id4_0_rdata = ram_w32_l4096_id4_0_rdata_out;
  reg [32-1:0] ram_w32_l4096_id4_1_rdata_out;
  assign ram_w32_l4096_id4_1_rdata = ram_w32_l4096_id4_1_rdata_out;
  reg [32-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w32_l4096_id4_0_enable) begin
      if(ram_w32_l4096_id4_0_wenable) begin
        mem[ram_w32_l4096_id4_0_addr] <= ram_w32_l4096_id4_0_wdata;
        ram_w32_l4096_id4_0_rdata_out <= ram_w32_l4096_id4_0_wdata;
      end else begin
        ram_w32_l4096_id4_0_rdata_out <= mem[ram_w32_l4096_id4_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l4096_id4_1_enable) begin
      if(ram_w32_l4096_id4_1_wenable) begin
        mem[ram_w32_l4096_id4_1_addr] <= ram_w32_l4096_id4_1_wdata;
        ram_w32_l4096_id4_1_rdata_out <= ram_w32_l4096_id4_1_wdata;
      end else begin
        ram_w32_l4096_id4_1_rdata_out <= mem[ram_w32_l4096_id4_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l4096_id5
(
  input CLK,
  input [12-1:0] ram_w32_l4096_id5_0_addr,
  output [32-1:0] ram_w32_l4096_id5_0_rdata,
  input [32-1:0] ram_w32_l4096_id5_0_wdata,
  input ram_w32_l4096_id5_0_wenable,
  input ram_w32_l4096_id5_0_enable,
  input [12-1:0] ram_w32_l4096_id5_1_addr,
  output [32-1:0] ram_w32_l4096_id5_1_rdata,
  input [32-1:0] ram_w32_l4096_id5_1_wdata,
  input ram_w32_l4096_id5_1_wenable,
  input ram_w32_l4096_id5_1_enable
);

  reg [32-1:0] ram_w32_l4096_id5_0_rdata_out;
  assign ram_w32_l4096_id5_0_rdata = ram_w32_l4096_id5_0_rdata_out;
  reg [32-1:0] ram_w32_l4096_id5_1_rdata_out;
  assign ram_w32_l4096_id5_1_rdata = ram_w32_l4096_id5_1_rdata_out;
  reg [32-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w32_l4096_id5_0_enable) begin
      if(ram_w32_l4096_id5_0_wenable) begin
        mem[ram_w32_l4096_id5_0_addr] <= ram_w32_l4096_id5_0_wdata;
        ram_w32_l4096_id5_0_rdata_out <= ram_w32_l4096_id5_0_wdata;
      end else begin
        ram_w32_l4096_id5_0_rdata_out <= mem[ram_w32_l4096_id5_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l4096_id5_1_enable) begin
      if(ram_w32_l4096_id5_1_wenable) begin
        mem[ram_w32_l4096_id5_1_addr] <= ram_w32_l4096_id5_1_wdata;
        ram_w32_l4096_id5_1_rdata_out <= ram_w32_l4096_id5_1_wdata;
      end else begin
        ram_w32_l4096_id5_1_rdata_out <= mem[ram_w32_l4096_id5_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l4096_id6
(
  input CLK,
  input [12-1:0] ram_w32_l4096_id6_0_addr,
  output [32-1:0] ram_w32_l4096_id6_0_rdata,
  input [32-1:0] ram_w32_l4096_id6_0_wdata,
  input ram_w32_l4096_id6_0_wenable,
  input ram_w32_l4096_id6_0_enable,
  input [12-1:0] ram_w32_l4096_id6_1_addr,
  output [32-1:0] ram_w32_l4096_id6_1_rdata,
  input [32-1:0] ram_w32_l4096_id6_1_wdata,
  input ram_w32_l4096_id6_1_wenable,
  input ram_w32_l4096_id6_1_enable
);

  reg [32-1:0] ram_w32_l4096_id6_0_rdata_out;
  assign ram_w32_l4096_id6_0_rdata = ram_w32_l4096_id6_0_rdata_out;
  reg [32-1:0] ram_w32_l4096_id6_1_rdata_out;
  assign ram_w32_l4096_id6_1_rdata = ram_w32_l4096_id6_1_rdata_out;
  reg [32-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w32_l4096_id6_0_enable) begin
      if(ram_w32_l4096_id6_0_wenable) begin
        mem[ram_w32_l4096_id6_0_addr] <= ram_w32_l4096_id6_0_wdata;
        ram_w32_l4096_id6_0_rdata_out <= ram_w32_l4096_id6_0_wdata;
      end else begin
        ram_w32_l4096_id6_0_rdata_out <= mem[ram_w32_l4096_id6_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l4096_id6_1_enable) begin
      if(ram_w32_l4096_id6_1_wenable) begin
        mem[ram_w32_l4096_id6_1_addr] <= ram_w32_l4096_id6_1_wdata;
        ram_w32_l4096_id6_1_rdata_out <= ram_w32_l4096_id6_1_wdata;
      end else begin
        ram_w32_l4096_id6_1_rdata_out <= mem[ram_w32_l4096_id6_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l4096_id7
(
  input CLK,
  input [12-1:0] ram_w32_l4096_id7_0_addr,
  output [32-1:0] ram_w32_l4096_id7_0_rdata,
  input [32-1:0] ram_w32_l4096_id7_0_wdata,
  input ram_w32_l4096_id7_0_wenable,
  input ram_w32_l4096_id7_0_enable,
  input [12-1:0] ram_w32_l4096_id7_1_addr,
  output [32-1:0] ram_w32_l4096_id7_1_rdata,
  input [32-1:0] ram_w32_l4096_id7_1_wdata,
  input ram_w32_l4096_id7_1_wenable,
  input ram_w32_l4096_id7_1_enable
);

  reg [32-1:0] ram_w32_l4096_id7_0_rdata_out;
  assign ram_w32_l4096_id7_0_rdata = ram_w32_l4096_id7_0_rdata_out;
  reg [32-1:0] ram_w32_l4096_id7_1_rdata_out;
  assign ram_w32_l4096_id7_1_rdata = ram_w32_l4096_id7_1_rdata_out;
  reg [32-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w32_l4096_id7_0_enable) begin
      if(ram_w32_l4096_id7_0_wenable) begin
        mem[ram_w32_l4096_id7_0_addr] <= ram_w32_l4096_id7_0_wdata;
        ram_w32_l4096_id7_0_rdata_out <= ram_w32_l4096_id7_0_wdata;
      end else begin
        ram_w32_l4096_id7_0_rdata_out <= mem[ram_w32_l4096_id7_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l4096_id7_1_enable) begin
      if(ram_w32_l4096_id7_1_wenable) begin
        mem[ram_w32_l4096_id7_1_addr] <= ram_w32_l4096_id7_1_wdata;
        ram_w32_l4096_id7_1_rdata_out <= ram_w32_l4096_id7_1_wdata;
      end else begin
        ram_w32_l4096_id7_1_rdata_out <= mem[ram_w32_l4096_id7_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l4096_id8
(
  input CLK,
  input [12-1:0] ram_w32_l4096_id8_0_addr,
  output [32-1:0] ram_w32_l4096_id8_0_rdata,
  input [32-1:0] ram_w32_l4096_id8_0_wdata,
  input ram_w32_l4096_id8_0_wenable,
  input ram_w32_l4096_id8_0_enable,
  input [12-1:0] ram_w32_l4096_id8_1_addr,
  output [32-1:0] ram_w32_l4096_id8_1_rdata,
  input [32-1:0] ram_w32_l4096_id8_1_wdata,
  input ram_w32_l4096_id8_1_wenable,
  input ram_w32_l4096_id8_1_enable
);

  reg [32-1:0] ram_w32_l4096_id8_0_rdata_out;
  assign ram_w32_l4096_id8_0_rdata = ram_w32_l4096_id8_0_rdata_out;
  reg [32-1:0] ram_w32_l4096_id8_1_rdata_out;
  assign ram_w32_l4096_id8_1_rdata = ram_w32_l4096_id8_1_rdata_out;
  reg [32-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w32_l4096_id8_0_enable) begin
      if(ram_w32_l4096_id8_0_wenable) begin
        mem[ram_w32_l4096_id8_0_addr] <= ram_w32_l4096_id8_0_wdata;
        ram_w32_l4096_id8_0_rdata_out <= ram_w32_l4096_id8_0_wdata;
      end else begin
        ram_w32_l4096_id8_0_rdata_out <= mem[ram_w32_l4096_id8_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l4096_id8_1_enable) begin
      if(ram_w32_l4096_id8_1_wenable) begin
        mem[ram_w32_l4096_id8_1_addr] <= ram_w32_l4096_id8_1_wdata;
        ram_w32_l4096_id8_1_rdata_out <= ram_w32_l4096_id8_1_wdata;
      end else begin
        ram_w32_l4096_id8_1_rdata_out <= mem[ram_w32_l4096_id8_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l1024_id0
(
  input CLK,
  input [10-1:0] ram_w32_l1024_id0_0_addr,
  output [32-1:0] ram_w32_l1024_id0_0_rdata,
  input [32-1:0] ram_w32_l1024_id0_0_wdata,
  input ram_w32_l1024_id0_0_wenable,
  input ram_w32_l1024_id0_0_enable,
  input [10-1:0] ram_w32_l1024_id0_1_addr,
  output [32-1:0] ram_w32_l1024_id0_1_rdata,
  input [32-1:0] ram_w32_l1024_id0_1_wdata,
  input ram_w32_l1024_id0_1_wenable,
  input ram_w32_l1024_id0_1_enable
);

  reg [32-1:0] ram_w32_l1024_id0_0_rdata_out;
  assign ram_w32_l1024_id0_0_rdata = ram_w32_l1024_id0_0_rdata_out;
  reg [32-1:0] ram_w32_l1024_id0_1_rdata_out;
  assign ram_w32_l1024_id0_1_rdata = ram_w32_l1024_id0_1_rdata_out;
  reg [32-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w32_l1024_id0_0_enable) begin
      if(ram_w32_l1024_id0_0_wenable) begin
        mem[ram_w32_l1024_id0_0_addr] <= ram_w32_l1024_id0_0_wdata;
        ram_w32_l1024_id0_0_rdata_out <= ram_w32_l1024_id0_0_wdata;
      end else begin
        ram_w32_l1024_id0_0_rdata_out <= mem[ram_w32_l1024_id0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l1024_id0_1_enable) begin
      if(ram_w32_l1024_id0_1_wenable) begin
        mem[ram_w32_l1024_id0_1_addr] <= ram_w32_l1024_id0_1_wdata;
        ram_w32_l1024_id0_1_rdata_out <= ram_w32_l1024_id0_1_wdata;
      end else begin
        ram_w32_l1024_id0_1_rdata_out <= mem[ram_w32_l1024_id0_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l1024_id1
(
  input CLK,
  input [10-1:0] ram_w32_l1024_id1_0_addr,
  output [32-1:0] ram_w32_l1024_id1_0_rdata,
  input [32-1:0] ram_w32_l1024_id1_0_wdata,
  input ram_w32_l1024_id1_0_wenable,
  input ram_w32_l1024_id1_0_enable,
  input [10-1:0] ram_w32_l1024_id1_1_addr,
  output [32-1:0] ram_w32_l1024_id1_1_rdata,
  input [32-1:0] ram_w32_l1024_id1_1_wdata,
  input ram_w32_l1024_id1_1_wenable,
  input ram_w32_l1024_id1_1_enable
);

  reg [32-1:0] ram_w32_l1024_id1_0_rdata_out;
  assign ram_w32_l1024_id1_0_rdata = ram_w32_l1024_id1_0_rdata_out;
  reg [32-1:0] ram_w32_l1024_id1_1_rdata_out;
  assign ram_w32_l1024_id1_1_rdata = ram_w32_l1024_id1_1_rdata_out;
  reg [32-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w32_l1024_id1_0_enable) begin
      if(ram_w32_l1024_id1_0_wenable) begin
        mem[ram_w32_l1024_id1_0_addr] <= ram_w32_l1024_id1_0_wdata;
        ram_w32_l1024_id1_0_rdata_out <= ram_w32_l1024_id1_0_wdata;
      end else begin
        ram_w32_l1024_id1_0_rdata_out <= mem[ram_w32_l1024_id1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l1024_id1_1_enable) begin
      if(ram_w32_l1024_id1_1_wenable) begin
        mem[ram_w32_l1024_id1_1_addr] <= ram_w32_l1024_id1_1_wdata;
        ram_w32_l1024_id1_1_rdata_out <= ram_w32_l1024_id1_1_wdata;
      end else begin
        ram_w32_l1024_id1_1_rdata_out <= mem[ram_w32_l1024_id1_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l1024_id2
(
  input CLK,
  input [10-1:0] ram_w32_l1024_id2_0_addr,
  output [32-1:0] ram_w32_l1024_id2_0_rdata,
  input [32-1:0] ram_w32_l1024_id2_0_wdata,
  input ram_w32_l1024_id2_0_wenable,
  input ram_w32_l1024_id2_0_enable,
  input [10-1:0] ram_w32_l1024_id2_1_addr,
  output [32-1:0] ram_w32_l1024_id2_1_rdata,
  input [32-1:0] ram_w32_l1024_id2_1_wdata,
  input ram_w32_l1024_id2_1_wenable,
  input ram_w32_l1024_id2_1_enable
);

  reg [32-1:0] ram_w32_l1024_id2_0_rdata_out;
  assign ram_w32_l1024_id2_0_rdata = ram_w32_l1024_id2_0_rdata_out;
  reg [32-1:0] ram_w32_l1024_id2_1_rdata_out;
  assign ram_w32_l1024_id2_1_rdata = ram_w32_l1024_id2_1_rdata_out;
  reg [32-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w32_l1024_id2_0_enable) begin
      if(ram_w32_l1024_id2_0_wenable) begin
        mem[ram_w32_l1024_id2_0_addr] <= ram_w32_l1024_id2_0_wdata;
        ram_w32_l1024_id2_0_rdata_out <= ram_w32_l1024_id2_0_wdata;
      end else begin
        ram_w32_l1024_id2_0_rdata_out <= mem[ram_w32_l1024_id2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l1024_id2_1_enable) begin
      if(ram_w32_l1024_id2_1_wenable) begin
        mem[ram_w32_l1024_id2_1_addr] <= ram_w32_l1024_id2_1_wdata;
        ram_w32_l1024_id2_1_rdata_out <= ram_w32_l1024_id2_1_wdata;
      end else begin
        ram_w32_l1024_id2_1_rdata_out <= mem[ram_w32_l1024_id2_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l1024_id3
(
  input CLK,
  input [10-1:0] ram_w32_l1024_id3_0_addr,
  output [32-1:0] ram_w32_l1024_id3_0_rdata,
  input [32-1:0] ram_w32_l1024_id3_0_wdata,
  input ram_w32_l1024_id3_0_wenable,
  input ram_w32_l1024_id3_0_enable,
  input [10-1:0] ram_w32_l1024_id3_1_addr,
  output [32-1:0] ram_w32_l1024_id3_1_rdata,
  input [32-1:0] ram_w32_l1024_id3_1_wdata,
  input ram_w32_l1024_id3_1_wenable,
  input ram_w32_l1024_id3_1_enable
);

  reg [32-1:0] ram_w32_l1024_id3_0_rdata_out;
  assign ram_w32_l1024_id3_0_rdata = ram_w32_l1024_id3_0_rdata_out;
  reg [32-1:0] ram_w32_l1024_id3_1_rdata_out;
  assign ram_w32_l1024_id3_1_rdata = ram_w32_l1024_id3_1_rdata_out;
  reg [32-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w32_l1024_id3_0_enable) begin
      if(ram_w32_l1024_id3_0_wenable) begin
        mem[ram_w32_l1024_id3_0_addr] <= ram_w32_l1024_id3_0_wdata;
        ram_w32_l1024_id3_0_rdata_out <= ram_w32_l1024_id3_0_wdata;
      end else begin
        ram_w32_l1024_id3_0_rdata_out <= mem[ram_w32_l1024_id3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l1024_id3_1_enable) begin
      if(ram_w32_l1024_id3_1_wenable) begin
        mem[ram_w32_l1024_id3_1_addr] <= ram_w32_l1024_id3_1_wdata;
        ram_w32_l1024_id3_1_rdata_out <= ram_w32_l1024_id3_1_wdata;
      end else begin
        ram_w32_l1024_id3_1_rdata_out <= mem[ram_w32_l1024_id3_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l1024_id4
(
  input CLK,
  input [10-1:0] ram_w32_l1024_id4_0_addr,
  output [32-1:0] ram_w32_l1024_id4_0_rdata,
  input [32-1:0] ram_w32_l1024_id4_0_wdata,
  input ram_w32_l1024_id4_0_wenable,
  input ram_w32_l1024_id4_0_enable,
  input [10-1:0] ram_w32_l1024_id4_1_addr,
  output [32-1:0] ram_w32_l1024_id4_1_rdata,
  input [32-1:0] ram_w32_l1024_id4_1_wdata,
  input ram_w32_l1024_id4_1_wenable,
  input ram_w32_l1024_id4_1_enable
);

  reg [32-1:0] ram_w32_l1024_id4_0_rdata_out;
  assign ram_w32_l1024_id4_0_rdata = ram_w32_l1024_id4_0_rdata_out;
  reg [32-1:0] ram_w32_l1024_id4_1_rdata_out;
  assign ram_w32_l1024_id4_1_rdata = ram_w32_l1024_id4_1_rdata_out;
  reg [32-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w32_l1024_id4_0_enable) begin
      if(ram_w32_l1024_id4_0_wenable) begin
        mem[ram_w32_l1024_id4_0_addr] <= ram_w32_l1024_id4_0_wdata;
        ram_w32_l1024_id4_0_rdata_out <= ram_w32_l1024_id4_0_wdata;
      end else begin
        ram_w32_l1024_id4_0_rdata_out <= mem[ram_w32_l1024_id4_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l1024_id4_1_enable) begin
      if(ram_w32_l1024_id4_1_wenable) begin
        mem[ram_w32_l1024_id4_1_addr] <= ram_w32_l1024_id4_1_wdata;
        ram_w32_l1024_id4_1_rdata_out <= ram_w32_l1024_id4_1_wdata;
      end else begin
        ram_w32_l1024_id4_1_rdata_out <= mem[ram_w32_l1024_id4_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l1024_id5
(
  input CLK,
  input [10-1:0] ram_w32_l1024_id5_0_addr,
  output [32-1:0] ram_w32_l1024_id5_0_rdata,
  input [32-1:0] ram_w32_l1024_id5_0_wdata,
  input ram_w32_l1024_id5_0_wenable,
  input ram_w32_l1024_id5_0_enable,
  input [10-1:0] ram_w32_l1024_id5_1_addr,
  output [32-1:0] ram_w32_l1024_id5_1_rdata,
  input [32-1:0] ram_w32_l1024_id5_1_wdata,
  input ram_w32_l1024_id5_1_wenable,
  input ram_w32_l1024_id5_1_enable
);

  reg [32-1:0] ram_w32_l1024_id5_0_rdata_out;
  assign ram_w32_l1024_id5_0_rdata = ram_w32_l1024_id5_0_rdata_out;
  reg [32-1:0] ram_w32_l1024_id5_1_rdata_out;
  assign ram_w32_l1024_id5_1_rdata = ram_w32_l1024_id5_1_rdata_out;
  reg [32-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w32_l1024_id5_0_enable) begin
      if(ram_w32_l1024_id5_0_wenable) begin
        mem[ram_w32_l1024_id5_0_addr] <= ram_w32_l1024_id5_0_wdata;
        ram_w32_l1024_id5_0_rdata_out <= ram_w32_l1024_id5_0_wdata;
      end else begin
        ram_w32_l1024_id5_0_rdata_out <= mem[ram_w32_l1024_id5_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l1024_id5_1_enable) begin
      if(ram_w32_l1024_id5_1_wenable) begin
        mem[ram_w32_l1024_id5_1_addr] <= ram_w32_l1024_id5_1_wdata;
        ram_w32_l1024_id5_1_rdata_out <= ram_w32_l1024_id5_1_wdata;
      end else begin
        ram_w32_l1024_id5_1_rdata_out <= mem[ram_w32_l1024_id5_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l1024_id6
(
  input CLK,
  input [10-1:0] ram_w32_l1024_id6_0_addr,
  output [32-1:0] ram_w32_l1024_id6_0_rdata,
  input [32-1:0] ram_w32_l1024_id6_0_wdata,
  input ram_w32_l1024_id6_0_wenable,
  input ram_w32_l1024_id6_0_enable,
  input [10-1:0] ram_w32_l1024_id6_1_addr,
  output [32-1:0] ram_w32_l1024_id6_1_rdata,
  input [32-1:0] ram_w32_l1024_id6_1_wdata,
  input ram_w32_l1024_id6_1_wenable,
  input ram_w32_l1024_id6_1_enable
);

  reg [32-1:0] ram_w32_l1024_id6_0_rdata_out;
  assign ram_w32_l1024_id6_0_rdata = ram_w32_l1024_id6_0_rdata_out;
  reg [32-1:0] ram_w32_l1024_id6_1_rdata_out;
  assign ram_w32_l1024_id6_1_rdata = ram_w32_l1024_id6_1_rdata_out;
  reg [32-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w32_l1024_id6_0_enable) begin
      if(ram_w32_l1024_id6_0_wenable) begin
        mem[ram_w32_l1024_id6_0_addr] <= ram_w32_l1024_id6_0_wdata;
        ram_w32_l1024_id6_0_rdata_out <= ram_w32_l1024_id6_0_wdata;
      end else begin
        ram_w32_l1024_id6_0_rdata_out <= mem[ram_w32_l1024_id6_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l1024_id6_1_enable) begin
      if(ram_w32_l1024_id6_1_wenable) begin
        mem[ram_w32_l1024_id6_1_addr] <= ram_w32_l1024_id6_1_wdata;
        ram_w32_l1024_id6_1_rdata_out <= ram_w32_l1024_id6_1_wdata;
      end else begin
        ram_w32_l1024_id6_1_rdata_out <= mem[ram_w32_l1024_id6_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l1024_id7
(
  input CLK,
  input [10-1:0] ram_w32_l1024_id7_0_addr,
  output [32-1:0] ram_w32_l1024_id7_0_rdata,
  input [32-1:0] ram_w32_l1024_id7_0_wdata,
  input ram_w32_l1024_id7_0_wenable,
  input ram_w32_l1024_id7_0_enable,
  input [10-1:0] ram_w32_l1024_id7_1_addr,
  output [32-1:0] ram_w32_l1024_id7_1_rdata,
  input [32-1:0] ram_w32_l1024_id7_1_wdata,
  input ram_w32_l1024_id7_1_wenable,
  input ram_w32_l1024_id7_1_enable
);

  reg [32-1:0] ram_w32_l1024_id7_0_rdata_out;
  assign ram_w32_l1024_id7_0_rdata = ram_w32_l1024_id7_0_rdata_out;
  reg [32-1:0] ram_w32_l1024_id7_1_rdata_out;
  assign ram_w32_l1024_id7_1_rdata = ram_w32_l1024_id7_1_rdata_out;
  reg [32-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w32_l1024_id7_0_enable) begin
      if(ram_w32_l1024_id7_0_wenable) begin
        mem[ram_w32_l1024_id7_0_addr] <= ram_w32_l1024_id7_0_wdata;
        ram_w32_l1024_id7_0_rdata_out <= ram_w32_l1024_id7_0_wdata;
      end else begin
        ram_w32_l1024_id7_0_rdata_out <= mem[ram_w32_l1024_id7_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l1024_id7_1_enable) begin
      if(ram_w32_l1024_id7_1_wenable) begin
        mem[ram_w32_l1024_id7_1_addr] <= ram_w32_l1024_id7_1_wdata;
        ram_w32_l1024_id7_1_rdata_out <= ram_w32_l1024_id7_1_wdata;
      end else begin
        ram_w32_l1024_id7_1_rdata_out <= mem[ram_w32_l1024_id7_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l1024_id8
(
  input CLK,
  input [10-1:0] ram_w32_l1024_id8_0_addr,
  output [32-1:0] ram_w32_l1024_id8_0_rdata,
  input [32-1:0] ram_w32_l1024_id8_0_wdata,
  input ram_w32_l1024_id8_0_wenable,
  input ram_w32_l1024_id8_0_enable,
  input [10-1:0] ram_w32_l1024_id8_1_addr,
  output [32-1:0] ram_w32_l1024_id8_1_rdata,
  input [32-1:0] ram_w32_l1024_id8_1_wdata,
  input ram_w32_l1024_id8_1_wenable,
  input ram_w32_l1024_id8_1_enable
);

  reg [32-1:0] ram_w32_l1024_id8_0_rdata_out;
  assign ram_w32_l1024_id8_0_rdata = ram_w32_l1024_id8_0_rdata_out;
  reg [32-1:0] ram_w32_l1024_id8_1_rdata_out;
  assign ram_w32_l1024_id8_1_rdata = ram_w32_l1024_id8_1_rdata_out;
  reg [32-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w32_l1024_id8_0_enable) begin
      if(ram_w32_l1024_id8_0_wenable) begin
        mem[ram_w32_l1024_id8_0_addr] <= ram_w32_l1024_id8_0_wdata;
        ram_w32_l1024_id8_0_rdata_out <= ram_w32_l1024_id8_0_wdata;
      end else begin
        ram_w32_l1024_id8_0_rdata_out <= mem[ram_w32_l1024_id8_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l1024_id8_1_enable) begin
      if(ram_w32_l1024_id8_1_wenable) begin
        mem[ram_w32_l1024_id8_1_addr] <= ram_w32_l1024_id8_1_wdata;
        ram_w32_l1024_id8_1_rdata_out <= ram_w32_l1024_id8_1_wdata;
      end else begin
        ram_w32_l1024_id8_1_rdata_out <= mem[ram_w32_l1024_id8_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l1024_id9
(
  input CLK,
  input [10-1:0] ram_w32_l1024_id9_0_addr,
  output [32-1:0] ram_w32_l1024_id9_0_rdata,
  input [32-1:0] ram_w32_l1024_id9_0_wdata,
  input ram_w32_l1024_id9_0_wenable,
  input ram_w32_l1024_id9_0_enable,
  input [10-1:0] ram_w32_l1024_id9_1_addr,
  output [32-1:0] ram_w32_l1024_id9_1_rdata,
  input [32-1:0] ram_w32_l1024_id9_1_wdata,
  input ram_w32_l1024_id9_1_wenable,
  input ram_w32_l1024_id9_1_enable
);

  reg [32-1:0] ram_w32_l1024_id9_0_rdata_out;
  assign ram_w32_l1024_id9_0_rdata = ram_w32_l1024_id9_0_rdata_out;
  reg [32-1:0] ram_w32_l1024_id9_1_rdata_out;
  assign ram_w32_l1024_id9_1_rdata = ram_w32_l1024_id9_1_rdata_out;
  reg [32-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w32_l1024_id9_0_enable) begin
      if(ram_w32_l1024_id9_0_wenable) begin
        mem[ram_w32_l1024_id9_0_addr] <= ram_w32_l1024_id9_0_wdata;
        ram_w32_l1024_id9_0_rdata_out <= ram_w32_l1024_id9_0_wdata;
      end else begin
        ram_w32_l1024_id9_0_rdata_out <= mem[ram_w32_l1024_id9_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l1024_id9_1_enable) begin
      if(ram_w32_l1024_id9_1_wenable) begin
        mem[ram_w32_l1024_id9_1_addr] <= ram_w32_l1024_id9_1_wdata;
        ram_w32_l1024_id9_1_rdata_out <= ram_w32_l1024_id9_1_wdata;
      end else begin
        ram_w32_l1024_id9_1_rdata_out <= mem[ram_w32_l1024_id9_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l1024_id10
(
  input CLK,
  input [10-1:0] ram_w32_l1024_id10_0_addr,
  output [32-1:0] ram_w32_l1024_id10_0_rdata,
  input [32-1:0] ram_w32_l1024_id10_0_wdata,
  input ram_w32_l1024_id10_0_wenable,
  input ram_w32_l1024_id10_0_enable,
  input [10-1:0] ram_w32_l1024_id10_1_addr,
  output [32-1:0] ram_w32_l1024_id10_1_rdata,
  input [32-1:0] ram_w32_l1024_id10_1_wdata,
  input ram_w32_l1024_id10_1_wenable,
  input ram_w32_l1024_id10_1_enable
);

  reg [32-1:0] ram_w32_l1024_id10_0_rdata_out;
  assign ram_w32_l1024_id10_0_rdata = ram_w32_l1024_id10_0_rdata_out;
  reg [32-1:0] ram_w32_l1024_id10_1_rdata_out;
  assign ram_w32_l1024_id10_1_rdata = ram_w32_l1024_id10_1_rdata_out;
  reg [32-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w32_l1024_id10_0_enable) begin
      if(ram_w32_l1024_id10_0_wenable) begin
        mem[ram_w32_l1024_id10_0_addr] <= ram_w32_l1024_id10_0_wdata;
        ram_w32_l1024_id10_0_rdata_out <= ram_w32_l1024_id10_0_wdata;
      end else begin
        ram_w32_l1024_id10_0_rdata_out <= mem[ram_w32_l1024_id10_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l1024_id10_1_enable) begin
      if(ram_w32_l1024_id10_1_wenable) begin
        mem[ram_w32_l1024_id10_1_addr] <= ram_w32_l1024_id10_1_wdata;
        ram_w32_l1024_id10_1_rdata_out <= ram_w32_l1024_id10_1_wdata;
      end else begin
        ram_w32_l1024_id10_1_rdata_out <= mem[ram_w32_l1024_id10_1_addr];
      end
    end 
  end


endmodule



module madd_0
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_0
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_0
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_1
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_1
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_1
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_2
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_2
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_2
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_3
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_3
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_3
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_4
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_4
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_4
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_5
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_5
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_5
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_6
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_6
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_6
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_7
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_7
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_7
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_8
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);


  madd_core_8
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_8
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [32-1:0] b,
  input [32-1:0] c,
  output [64-1:0] d
);

  reg signed [32-1:0] _a;
  reg signed [32-1:0] _b;
  reg signed [32-1:0] _c;
  wire signed [64-1:0] _mul;
  wire signed [64-1:0] _madd;
  reg signed [64-1:0] _pipe_madd0;
  reg signed [64-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module multiplier_0
(
  input CLK,
  input update,
  input [128-1:0] a,
  input [32-1:0] b,
  output [160-1:0] c
);


  multiplier_core_0
  mult
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c)
  );


endmodule



module multiplier_core_0
(
  input CLK,
  input update,
  input [128-1:0] a,
  input [32-1:0] b,
  output [160-1:0] c
);

  reg signed [128-1:0] _a;
  reg signed [32-1:0] _b;
  wire signed [160-1:0] _mul;
  reg signed [160-1:0] _pipe_mul0;
  reg signed [160-1:0] _pipe_mul1;
  assign _mul = _a * _b;
  assign c = _pipe_mul1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _pipe_mul0 <= _mul;
      _pipe_mul1 <= _pipe_mul0;
    end 
  end


endmodule



module multiplier_1
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [29-1:0] b,
  output [61-1:0] c
);


  multiplier_core_1
  mult
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c)
  );


endmodule



module multiplier_core_1
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [29-1:0] b,
  output [61-1:0] c
);

  reg signed [32-1:0] _a;
  reg signed [29-1:0] _b;
  wire signed [61-1:0] _mul;
  reg signed [61-1:0] _pipe_mul0;
  assign _mul = _a * _b;
  assign c = _pipe_mul0;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _pipe_mul0 <= _mul;
    end 
  end


endmodule

